/*
Computer Architecture Lab 4 - 22-01-2018
	Assignment : Full Associative Cache
					Byte addressable Cache with Full Associative mapping to the Memory
					Physical Address of 12 bits (2^12 Bytes) in Main Memory
									Width	x	Depth
					Memory Size	: 2^4 Byte	x	2^8 Lines
					Cache Size	: 2^4 Byte	x	2^4 Cache Blocks

	Module : Associative Mapped Cache
		-- Eshita Arza	(COE15B013)
		-- Akshay Kumar	(CED15I031)
*/

module associative_cache(addr, clk, enable, line, chk_hit, ByTe);

	input [11:0]addr;
	input clk;
	input enable;

	output reg[127:0]line;
	output [7:0]ByTe;
	output reg chk_hit;

	reg [127:0]mem_line[255:0]; //main memory
	reg [127:0]cache_line[15:0]; //cache memory
	reg [7:0]tag_array[15:0]; //tag array
	//reg [3:0]cache_blk; //mentions the specific cache block
	reg [7:0]random; //randomly generates a 8 bit address
	reg [7:0]temp; //stores the current mapping address value generated by random
	wire [15:0]hit;	

	wire [7:0]tag_inp; 
	wire [3:0]Block_Offset; 

	integer i, j;
	integer rand;

	always@ (enable)
	begin
		for(i = 0; i < 256; ++i)
			mem_line[i] = i;
	end

	always@(enable)
	begin
		rand = 256;
		for(j = 0; j < 16; ++j)
		begin
			random = $random(rand);
			tag_array[j][7:0] = random[7:0];
			temp[7:0] = random[7:0];
			cache_line[j] = mem_line[temp]; //storing main memeory data of address pointed by temp into cache at location j 
		end
	end

	assign tag_inp[7:0] = addr[11:4]; //assigning tag_inp value from input address
	assign Block_Offset[3:0] = addr[3:0];  //assigning Block_Offset value from input address

	comparator_a c0(tag_inp, tag_array[0], hit[0]);
	comparator_a c1(tag_inp, tag_array[1], hit[1]);
	comparator_a c2(tag_inp, tag_array[2], hit[2]);
	comparator_a c3(tag_inp, tag_array[3], hit[3]);
	comparator_a c4(tag_inp, tag_array[4], hit[4]);
	comparator_a c5(tag_inp, tag_array[5], hit[5]);
	comparator_a c6(tag_inp, tag_array[6], hit[6]);
	comparator_a c7(tag_inp, tag_array[7], hit[7]);
	comparator_a c8(tag_inp, tag_array[8], hit[8]);
	comparator_a c9(tag_inp, tag_array[9], hit[9]);
	comparator_a c10(tag_inp, tag_array[10], hit[10]);
	comparator_a c11(tag_inp, tag_array[11], hit[11]);
	comparator_a c12(tag_inp, tag_array[12], hit[12]);
	comparator_a c13(tag_inp, tag_array[13], hit[13]);
	comparator_a c14(tag_inp, tag_array[14], hit[14]);
	comparator_a c15(tag_inp, tag_array[15], hit[15]);

	always@(negedge clk)
	begin
		chk_hit = hit[0] | hit[1] | hit[2] | hit[3] | hit[4] | hit[5] | hit[6] | hit[7] | hit[8] | hit[9] | hit[10] | hit[11] | hit[12] | hit[13] | hit[14] | hit[15];

		if(chk_hit == 1'b1)
		begin
			if(hit[0] == 1'b1)
			 	line[127:0] = cache_line[0][127:0];
			
			else if(hit[1] == 1'b1)
			 	line[127:0] = cache_line[1][127:0];
			
			else if(hit[2] == 1'b1)
			 	line[127:0] = cache_line[2][127:0];
			
			else if(hit[3] == 1'b1)
			 	line[127:0] = cache_line[3][127:0];
			
			else if(hit[4] == 1'b1)
			 	line[127:0] = cache_line[4][127:0];
			
			else if(hit[5] == 1'b1)
			 	line[127:0] = cache_line[5][127:0];
			
			else if(hit[6] == 1'b1)
			 	line[127:0] = cache_line[6][127:0];
			
			else if(hit[7] == 1'b1)
			 	line[127:0] = cache_line[7][127:0];
			
			else if(hit[8] == 1'b1)
			 	line[127:0] = cache_line[8][127:0];
			
			else if(hit[9] == 1'b1)
			 	line[127:0] = cache_line[9][127:0];
			
			else if(hit[10] == 1'b1)
			 	line[127:0] = cache_line[10][127:0];
			
			else if(hit[11] == 1'b1)
			 	line[127:0] = cache_line[11][127:0];
			
			else if(hit[12] == 1'b1)
			 	line[127:0] = cache_line[12][127:0];
			
			else if(hit[13] == 1'b1)
			 	line[127:0] = cache_line[13][127:0];
			
			else if(hit[14] == 1'b1)
			 	line[127:0] = cache_line[14][127:0];
			
			else if(hit[15] == 1'b1)
			 	line[127:0] = cache_line[15][127:0];
		end
		
		else if(chk_hit == 1'b0)
		begin
			rand = 16;
			random = $random(rand);
			j = random;
			tag_array[j][7:0] = tag_inp[7:0];
			cache_line[j][127:0] = mem_line[tag_inp[7:0]];
			line[127:0] = cache_line[j][127:0];	
		end
	end

	Offset_2_Byte b(line, Block_Offset, ByTe);

endmodule // associative_cache