/*
Computer Architecture Lab 3 - 15-01-2018
	Assignment : Direct Mapped Cache
					Byte addressable Cache with direct mapping to the Memory
					Physical Address of 32 bits (2^32 Bytes) in Main Memory
									Width	x	Depth
					Memory Size	: 2^8 Byte	x	2^24 Lines
					Cache Size	: 2^8 Byte	x	2^8 Cache Blocks
					Cache to Memory Mapping Ratio : 1 : 2^16

	Module : Direct Mapped Cache
		-- Eshita Arza	(COE15B013)
		-- Akshay Kumar	(CED15I031)
*/

module direct_cache(clk, addr, enable, line, hit, ByTe);

	input [31:0]addr;
	input clk;
	input enable;

	output reg [2047:0]line;
	output hit;
	output [7:0]ByTe;
	// reg [7:0]linterest;
	//output [7:0]loi;

	reg [2047:0]mem_line[16777215:0];
	reg [2047:0]cache_line[255:0];
	reg [15:0]tag_array[255:0];
	reg [7:0]temp_line;
	reg [23:0]map_line[255:0];
	reg [15:0]random;
	reg [7:0]cache_blk;

	wire chk;
	wire [23:0]line_addr;
	wire [7:0]line_interest;
	wire [15:0]tag_inp;
	wire [7:0]Block_Offset;

	integer i, j, k, rand, temp, flag;

	assign chk = 1'b0;
	always@ (enable)
	begin
		for(i = 0; i < 16777216; i = i + 1)
			mem_line[i] = i;
		//flag = 1;
	end

	always@ (enable)
	begin
		rand = 65536;
		for(j = 0; j < 256; j = j + 1)
		begin
			random = $random(rand);
			cache_blk = j;
			map_line[j][7:0] = cache_blk[7:0];
			map_line[j][23:8] = random[15:0];
			tag_array[j][15:0] = map_line[j][23:8];
			temp = map_line[j];
			cache_line[j] = mem_line[temp];
		end
	end

	/* extracting values of interest for the search from the address input */
	assign line_addr[23:0] = addr[31:8];
	assign tag_inp[15:0] = addr[31:16];
	assign line_interest[7:0] = addr[15:8];
	assign Block_Offset[7:0] = addr[7:0];

	//assign line_addr = addr[31:8];
	//assign tag_inp = addr[];

	//always@ (negedge clk) begin
	comparator c(tag_inp, tag_array[line_interest], hit, chk);

	/*always@(negedge clk)
	begin
	cache_line[0] = mem_line[0];
	line = cache_line[0];
	end*/
	//end

	//assign chk = 1'b1;

	/* in case of cache miss, load the respective line from Memory */
	always@ (negedge clk)
	begin
				k = line_interest;
		//if(chk == 1'b1)
		//	begin
				cache_line[k][0] = (mem_line[line_addr][0] & (~hit)) | (cache_line[k][0] & (hit));
				cache_line[k][1] = (mem_line[line_addr][1] & (~hit)) | (cache_line[k][1] & (hit));
				cache_line[k][2] = (mem_line[line_addr][2] & (~hit)) | (cache_line[k][2] & (hit));
				cache_line[k][3] = (mem_line[line_addr][3] & (~hit)) | (cache_line[k][3] & (hit));
				cache_line[k][4] = (mem_line[line_addr][4] & (~hit)) | (cache_line[k][4] & (hit));
				cache_line[k][5] = (mem_line[line_addr][5] & (~hit)) | (cache_line[k][5] & (hit));
				cache_line[k][6] = (mem_line[line_addr][6] & (~hit)) | (cache_line[k][6] & (hit));
				cache_line[k][7] = (mem_line[line_addr][7] & (~hit)) | (cache_line[k][7] & (hit));
				cache_line[k][8] = (mem_line[line_addr][8] & (~hit)) | (cache_line[k][8] & (hit));
				cache_line[k][9] = (mem_line[line_addr][9] & (~hit)) | (cache_line[k][9] & (hit));
				cache_line[k][10] = (mem_line[line_addr][10] & (~hit)) | (cache_line[k][10] & (hit));
				cache_line[k][11] = (mem_line[line_addr][11] & (~hit)) | (cache_line[k][11] & (hit));
				cache_line[k][12] = (mem_line[line_addr][12] & (~hit)) | (cache_line[k][12] & (hit));
				cache_line[k][13] = (mem_line[line_addr][13] & (~hit)) | (cache_line[k][13] & (hit));
				cache_line[k][14] = (mem_line[line_addr][14] & (~hit)) | (cache_line[k][14] & (hit));
				cache_line[k][15] = (mem_line[line_addr][15] & (~hit)) | (cache_line[k][15] & (hit));
				cache_line[k][16] = (mem_line[line_addr][16] & (~hit)) | (cache_line[k][16] & (hit));
				cache_line[k][17] = (mem_line[line_addr][17] & (~hit)) | (cache_line[k][17] & (hit));
				cache_line[k][18] = (mem_line[line_addr][18] & (~hit)) | (cache_line[k][18] & (hit));
				cache_line[k][19] = (mem_line[line_addr][19] & (~hit)) | (cache_line[k][19] & (hit));
				cache_line[k][20] = (mem_line[line_addr][20] & (~hit)) | (cache_line[k][20] & (hit));
				cache_line[k][21] = (mem_line[line_addr][21] & (~hit)) | (cache_line[k][21] & (hit));
				cache_line[k][22] = (mem_line[line_addr][22] & (~hit)) | (cache_line[k][22] & (hit));
				cache_line[k][23] = (mem_line[line_addr][23] & (~hit)) | (cache_line[k][23] & (hit));
				cache_line[k][24] = (mem_line[line_addr][24] & (~hit)) | (cache_line[k][24] & (hit));
				cache_line[k][25] = (mem_line[line_addr][25] & (~hit)) | (cache_line[k][25] & (hit));
				cache_line[k][26] = (mem_line[line_addr][26] & (~hit)) | (cache_line[k][26] & (hit));
				cache_line[k][27] = (mem_line[line_addr][27] & (~hit)) | (cache_line[k][27] & (hit));
				cache_line[k][28] = (mem_line[line_addr][28] & (~hit)) | (cache_line[k][28] & (hit));
				cache_line[k][29] = (mem_line[line_addr][29] & (~hit)) | (cache_line[k][29] & (hit));
				cache_line[k][30] = (mem_line[line_addr][30] & (~hit)) | (cache_line[k][30] & (hit));
				cache_line[k][31] = (mem_line[line_addr][31] & (~hit)) | (cache_line[k][31] & (hit));
				cache_line[k][32] = (mem_line[line_addr][32] & (~hit)) | (cache_line[k][32] & (hit));
				cache_line[k][33] = (mem_line[line_addr][33] & (~hit)) | (cache_line[k][33] & (hit));
				cache_line[k][34] = (mem_line[line_addr][34] & (~hit)) | (cache_line[k][34] & (hit));
				cache_line[k][35] = (mem_line[line_addr][35] & (~hit)) | (cache_line[k][35] & (hit));
				cache_line[k][36] = (mem_line[line_addr][36] & (~hit)) | (cache_line[k][36] & (hit));
				cache_line[k][37] = (mem_line[line_addr][37] & (~hit)) | (cache_line[k][37] & (hit));
				cache_line[k][38] = (mem_line[line_addr][38] & (~hit)) | (cache_line[k][38] & (hit));
				cache_line[k][39] = (mem_line[line_addr][39] & (~hit)) | (cache_line[k][39] & (hit));
				cache_line[k][40] = (mem_line[line_addr][40] & (~hit)) | (cache_line[k][40] & (hit));
				cache_line[k][41] = (mem_line[line_addr][41] & (~hit)) | (cache_line[k][41] & (hit));
				cache_line[k][42] = (mem_line[line_addr][42] & (~hit)) | (cache_line[k][42] & (hit));
				cache_line[k][43] = (mem_line[line_addr][43] & (~hit)) | (cache_line[k][43] & (hit));
				cache_line[k][44] = (mem_line[line_addr][44] & (~hit)) | (cache_line[k][44] & (hit));
				cache_line[k][45] = (mem_line[line_addr][45] & (~hit)) | (cache_line[k][45] & (hit));
				cache_line[k][46] = (mem_line[line_addr][46] & (~hit)) | (cache_line[k][46] & (hit));
				cache_line[k][47] = (mem_line[line_addr][47] & (~hit)) | (cache_line[k][47] & (hit));
				cache_line[k][48] = (mem_line[line_addr][48] & (~hit)) | (cache_line[k][48] & (hit));
				cache_line[k][49] = (mem_line[line_addr][49] & (~hit)) | (cache_line[k][49] & (hit));
				cache_line[k][50] = (mem_line[line_addr][50] & (~hit)) | (cache_line[k][50] & (hit));
				cache_line[k][51] = (mem_line[line_addr][51] & (~hit)) | (cache_line[k][51] & (hit));
				cache_line[k][52] = (mem_line[line_addr][52] & (~hit)) | (cache_line[k][52] & (hit));
				cache_line[k][53] = (mem_line[line_addr][53] & (~hit)) | (cache_line[k][53] & (hit));
				cache_line[k][54] = (mem_line[line_addr][54] & (~hit)) | (cache_line[k][54] & (hit));
				cache_line[k][55] = (mem_line[line_addr][55] & (~hit)) | (cache_line[k][55] & (hit));
				cache_line[k][56] = (mem_line[line_addr][56] & (~hit)) | (cache_line[k][56] & (hit));
				cache_line[k][57] = (mem_line[line_addr][57] & (~hit)) | (cache_line[k][57] & (hit));
				cache_line[k][58] = (mem_line[line_addr][58] & (~hit)) | (cache_line[k][58] & (hit));
				cache_line[k][59] = (mem_line[line_addr][59] & (~hit)) | (cache_line[k][59] & (hit));
				cache_line[k][60] = (mem_line[line_addr][60] & (~hit)) | (cache_line[k][60] & (hit));
				cache_line[k][61] = (mem_line[line_addr][61] & (~hit)) | (cache_line[k][61] & (hit));
				cache_line[k][62] = (mem_line[line_addr][62] & (~hit)) | (cache_line[k][62] & (hit));
				cache_line[k][63] = (mem_line[line_addr][63] & (~hit)) | (cache_line[k][63] & (hit));
				cache_line[k][64] = (mem_line[line_addr][64] & (~hit)) | (cache_line[k][64] & (hit));
				cache_line[k][65] = (mem_line[line_addr][65] & (~hit)) | (cache_line[k][65] & (hit));
				cache_line[k][66] = (mem_line[line_addr][66] & (~hit)) | (cache_line[k][66] & (hit));
				cache_line[k][67] = (mem_line[line_addr][67] & (~hit)) | (cache_line[k][67] & (hit));
				cache_line[k][68] = (mem_line[line_addr][68] & (~hit)) | (cache_line[k][68] & (hit));
				cache_line[k][69] = (mem_line[line_addr][69] & (~hit)) | (cache_line[k][69] & (hit));
				cache_line[k][70] = (mem_line[line_addr][70] & (~hit)) | (cache_line[k][70] & (hit));
				cache_line[k][71] = (mem_line[line_addr][71] & (~hit)) | (cache_line[k][71] & (hit));
				cache_line[k][72] = (mem_line[line_addr][72] & (~hit)) | (cache_line[k][72] & (hit));
				cache_line[k][73] = (mem_line[line_addr][73] & (~hit)) | (cache_line[k][73] & (hit));
				cache_line[k][74] = (mem_line[line_addr][74] & (~hit)) | (cache_line[k][74] & (hit));
				cache_line[k][75] = (mem_line[line_addr][75] & (~hit)) | (cache_line[k][75] & (hit));
				cache_line[k][76] = (mem_line[line_addr][76] & (~hit)) | (cache_line[k][76] & (hit));
				cache_line[k][77] = (mem_line[line_addr][77] & (~hit)) | (cache_line[k][77] & (hit));
				cache_line[k][78] = (mem_line[line_addr][78] & (~hit)) | (cache_line[k][78] & (hit));
				cache_line[k][79] = (mem_line[line_addr][79] & (~hit)) | (cache_line[k][79] & (hit));
				cache_line[k][80] = (mem_line[line_addr][80] & (~hit)) | (cache_line[k][80] & (hit));
				cache_line[k][81] = (mem_line[line_addr][81] & (~hit)) | (cache_line[k][81] & (hit));
				cache_line[k][82] = (mem_line[line_addr][82] & (~hit)) | (cache_line[k][82] & (hit));
				cache_line[k][83] = (mem_line[line_addr][83] & (~hit)) | (cache_line[k][83] & (hit));
				cache_line[k][84] = (mem_line[line_addr][84] & (~hit)) | (cache_line[k][84] & (hit));
				cache_line[k][85] = (mem_line[line_addr][85] & (~hit)) | (cache_line[k][85] & (hit));
				cache_line[k][86] = (mem_line[line_addr][86] & (~hit)) | (cache_line[k][86] & (hit));
				cache_line[k][87] = (mem_line[line_addr][87] & (~hit)) | (cache_line[k][87] & (hit));
				cache_line[k][88] = (mem_line[line_addr][88] & (~hit)) | (cache_line[k][88] & (hit));
				cache_line[k][89] = (mem_line[line_addr][89] & (~hit)) | (cache_line[k][89] & (hit));
				cache_line[k][90] = (mem_line[line_addr][90] & (~hit)) | (cache_line[k][90] & (hit));
				cache_line[k][91] = (mem_line[line_addr][91] & (~hit)) | (cache_line[k][91] & (hit));
				cache_line[k][92] = (mem_line[line_addr][92] & (~hit)) | (cache_line[k][92] & (hit));
				cache_line[k][93] = (mem_line[line_addr][93] & (~hit)) | (cache_line[k][93] & (hit));
				cache_line[k][94] = (mem_line[line_addr][94] & (~hit)) | (cache_line[k][94] & (hit));
				cache_line[k][95] = (mem_line[line_addr][95] & (~hit)) | (cache_line[k][95] & (hit));
				cache_line[k][96] = (mem_line[line_addr][96] & (~hit)) | (cache_line[k][96] & (hit));
				cache_line[k][97] = (mem_line[line_addr][97] & (~hit)) | (cache_line[k][97] & (hit));
				cache_line[k][98] = (mem_line[line_addr][98] & (~hit)) | (cache_line[k][98] & (hit));
				cache_line[k][99] = (mem_line[line_addr][99] & (~hit)) | (cache_line[k][99] & (hit));
				cache_line[k][100] = (mem_line[line_addr][100] & (~hit)) | (cache_line[k][100] & (hit));
				cache_line[k][101] = (mem_line[line_addr][101] & (~hit)) | (cache_line[k][101] & (hit));
				cache_line[k][102] = (mem_line[line_addr][102] & (~hit)) | (cache_line[k][102] & (hit));
				cache_line[k][103] = (mem_line[line_addr][103] & (~hit)) | (cache_line[k][103] & (hit));
				cache_line[k][104] = (mem_line[line_addr][104] & (~hit)) | (cache_line[k][104] & (hit));
				cache_line[k][105] = (mem_line[line_addr][105] & (~hit)) | (cache_line[k][105] & (hit));
				cache_line[k][106] = (mem_line[line_addr][106] & (~hit)) | (cache_line[k][106] & (hit));
				cache_line[k][107] = (mem_line[line_addr][107] & (~hit)) | (cache_line[k][107] & (hit));
				cache_line[k][108] = (mem_line[line_addr][108] & (~hit)) | (cache_line[k][108] & (hit));
				cache_line[k][109] = (mem_line[line_addr][109] & (~hit)) | (cache_line[k][109] & (hit));
				cache_line[k][110] = (mem_line[line_addr][110] & (~hit)) | (cache_line[k][110] & (hit));
				cache_line[k][111] = (mem_line[line_addr][111] & (~hit)) | (cache_line[k][111] & (hit));
				cache_line[k][112] = (mem_line[line_addr][112] & (~hit)) | (cache_line[k][112] & (hit));
				cache_line[k][113] = (mem_line[line_addr][113] & (~hit)) | (cache_line[k][113] & (hit));
				cache_line[k][114] = (mem_line[line_addr][114] & (~hit)) | (cache_line[k][114] & (hit));
				cache_line[k][115] = (mem_line[line_addr][115] & (~hit)) | (cache_line[k][115] & (hit));
				cache_line[k][116] = (mem_line[line_addr][116] & (~hit)) | (cache_line[k][116] & (hit));
				cache_line[k][117] = (mem_line[line_addr][117] & (~hit)) | (cache_line[k][117] & (hit));
				cache_line[k][118] = (mem_line[line_addr][118] & (~hit)) | (cache_line[k][118] & (hit));
				cache_line[k][119] = (mem_line[line_addr][119] & (~hit)) | (cache_line[k][119] & (hit));
				cache_line[k][120] = (mem_line[line_addr][120] & (~hit)) | (cache_line[k][120] & (hit));
				cache_line[k][121] = (mem_line[line_addr][121] & (~hit)) | (cache_line[k][121] & (hit));
				cache_line[k][122] = (mem_line[line_addr][122] & (~hit)) | (cache_line[k][122] & (hit));
				cache_line[k][123] = (mem_line[line_addr][123] & (~hit)) | (cache_line[k][123] & (hit));
				cache_line[k][124] = (mem_line[line_addr][124] & (~hit)) | (cache_line[k][124] & (hit));
				cache_line[k][125] = (mem_line[line_addr][125] & (~hit)) | (cache_line[k][125] & (hit));
				cache_line[k][126] = (mem_line[line_addr][126] & (~hit)) | (cache_line[k][126] & (hit));
				cache_line[k][127] = (mem_line[line_addr][127] & (~hit)) | (cache_line[k][127] & (hit));
				cache_line[k][128] = (mem_line[line_addr][128] & (~hit)) | (cache_line[k][128] & (hit));
				cache_line[k][129] = (mem_line[line_addr][129] & (~hit)) | (cache_line[k][129] & (hit));
				cache_line[k][130] = (mem_line[line_addr][130] & (~hit)) | (cache_line[k][130] & (hit));
				cache_line[k][131] = (mem_line[line_addr][131] & (~hit)) | (cache_line[k][131] & (hit));
				cache_line[k][132] = (mem_line[line_addr][132] & (~hit)) | (cache_line[k][132] & (hit));
				cache_line[k][133] = (mem_line[line_addr][133] & (~hit)) | (cache_line[k][133] & (hit));
				cache_line[k][134] = (mem_line[line_addr][134] & (~hit)) | (cache_line[k][134] & (hit));
				cache_line[k][135] = (mem_line[line_addr][135] & (~hit)) | (cache_line[k][135] & (hit));
				cache_line[k][136] = (mem_line[line_addr][136] & (~hit)) | (cache_line[k][136] & (hit));
				cache_line[k][137] = (mem_line[line_addr][137] & (~hit)) | (cache_line[k][137] & (hit));
				cache_line[k][138] = (mem_line[line_addr][138] & (~hit)) | (cache_line[k][138] & (hit));
				cache_line[k][139] = (mem_line[line_addr][139] & (~hit)) | (cache_line[k][139] & (hit));
				cache_line[k][140] = (mem_line[line_addr][140] & (~hit)) | (cache_line[k][140] & (hit));
				cache_line[k][141] = (mem_line[line_addr][141] & (~hit)) | (cache_line[k][141] & (hit));
				cache_line[k][142] = (mem_line[line_addr][142] & (~hit)) | (cache_line[k][142] & (hit));
				cache_line[k][143] = (mem_line[line_addr][143] & (~hit)) | (cache_line[k][143] & (hit));
				cache_line[k][144] = (mem_line[line_addr][144] & (~hit)) | (cache_line[k][144] & (hit));
				cache_line[k][145] = (mem_line[line_addr][145] & (~hit)) | (cache_line[k][145] & (hit));
				cache_line[k][146] = (mem_line[line_addr][146] & (~hit)) | (cache_line[k][146] & (hit));
				cache_line[k][147] = (mem_line[line_addr][147] & (~hit)) | (cache_line[k][147] & (hit));
				cache_line[k][148] = (mem_line[line_addr][148] & (~hit)) | (cache_line[k][148] & (hit));
				cache_line[k][149] = (mem_line[line_addr][149] & (~hit)) | (cache_line[k][149] & (hit));
				cache_line[k][150] = (mem_line[line_addr][150] & (~hit)) | (cache_line[k][150] & (hit));
				cache_line[k][151] = (mem_line[line_addr][151] & (~hit)) | (cache_line[k][151] & (hit));
				cache_line[k][152] = (mem_line[line_addr][152] & (~hit)) | (cache_line[k][152] & (hit));
				cache_line[k][153] = (mem_line[line_addr][153] & (~hit)) | (cache_line[k][153] & (hit));
				cache_line[k][154] = (mem_line[line_addr][154] & (~hit)) | (cache_line[k][154] & (hit));
				cache_line[k][155] = (mem_line[line_addr][155] & (~hit)) | (cache_line[k][155] & (hit));
				cache_line[k][156] = (mem_line[line_addr][156] & (~hit)) | (cache_line[k][156] & (hit));
				cache_line[k][157] = (mem_line[line_addr][157] & (~hit)) | (cache_line[k][157] & (hit));
				cache_line[k][158] = (mem_line[line_addr][158] & (~hit)) | (cache_line[k][158] & (hit));
				cache_line[k][159] = (mem_line[line_addr][159] & (~hit)) | (cache_line[k][159] & (hit));
				cache_line[k][160] = (mem_line[line_addr][160] & (~hit)) | (cache_line[k][160] & (hit));
				cache_line[k][161] = (mem_line[line_addr][161] & (~hit)) | (cache_line[k][161] & (hit));
				cache_line[k][162] = (mem_line[line_addr][162] & (~hit)) | (cache_line[k][162] & (hit));
				cache_line[k][163] = (mem_line[line_addr][163] & (~hit)) | (cache_line[k][163] & (hit));
				cache_line[k][164] = (mem_line[line_addr][164] & (~hit)) | (cache_line[k][164] & (hit));
				cache_line[k][165] = (mem_line[line_addr][165] & (~hit)) | (cache_line[k][165] & (hit));
				cache_line[k][166] = (mem_line[line_addr][166] & (~hit)) | (cache_line[k][166] & (hit));
				cache_line[k][167] = (mem_line[line_addr][167] & (~hit)) | (cache_line[k][167] & (hit));
				cache_line[k][168] = (mem_line[line_addr][168] & (~hit)) | (cache_line[k][168] & (hit));
				cache_line[k][169] = (mem_line[line_addr][169] & (~hit)) | (cache_line[k][169] & (hit));
				cache_line[k][170] = (mem_line[line_addr][170] & (~hit)) | (cache_line[k][170] & (hit));
				cache_line[k][171] = (mem_line[line_addr][171] & (~hit)) | (cache_line[k][171] & (hit));
				cache_line[k][172] = (mem_line[line_addr][172] & (~hit)) | (cache_line[k][172] & (hit));
				cache_line[k][173] = (mem_line[line_addr][173] & (~hit)) | (cache_line[k][173] & (hit));
				cache_line[k][174] = (mem_line[line_addr][174] & (~hit)) | (cache_line[k][174] & (hit));
				cache_line[k][175] = (mem_line[line_addr][175] & (~hit)) | (cache_line[k][175] & (hit));
				cache_line[k][176] = (mem_line[line_addr][176] & (~hit)) | (cache_line[k][176] & (hit));
				cache_line[k][177] = (mem_line[line_addr][177] & (~hit)) | (cache_line[k][177] & (hit));
				cache_line[k][178] = (mem_line[line_addr][178] & (~hit)) | (cache_line[k][178] & (hit));
				cache_line[k][179] = (mem_line[line_addr][179] & (~hit)) | (cache_line[k][179] & (hit));
				cache_line[k][180] = (mem_line[line_addr][180] & (~hit)) | (cache_line[k][180] & (hit));
				cache_line[k][181] = (mem_line[line_addr][181] & (~hit)) | (cache_line[k][181] & (hit));
				cache_line[k][182] = (mem_line[line_addr][182] & (~hit)) | (cache_line[k][182] & (hit));
				cache_line[k][183] = (mem_line[line_addr][183] & (~hit)) | (cache_line[k][183] & (hit));
				cache_line[k][184] = (mem_line[line_addr][184] & (~hit)) | (cache_line[k][184] & (hit));
				cache_line[k][185] = (mem_line[line_addr][185] & (~hit)) | (cache_line[k][185] & (hit));
				cache_line[k][186] = (mem_line[line_addr][186] & (~hit)) | (cache_line[k][186] & (hit));
				cache_line[k][187] = (mem_line[line_addr][187] & (~hit)) | (cache_line[k][187] & (hit));
				cache_line[k][188] = (mem_line[line_addr][188] & (~hit)) | (cache_line[k][188] & (hit));
				cache_line[k][189] = (mem_line[line_addr][189] & (~hit)) | (cache_line[k][189] & (hit));
				cache_line[k][190] = (mem_line[line_addr][190] & (~hit)) | (cache_line[k][190] & (hit));
				cache_line[k][191] = (mem_line[line_addr][191] & (~hit)) | (cache_line[k][191] & (hit));
				cache_line[k][192] = (mem_line[line_addr][192] & (~hit)) | (cache_line[k][192] & (hit));
				cache_line[k][193] = (mem_line[line_addr][193] & (~hit)) | (cache_line[k][193] & (hit));
				cache_line[k][194] = (mem_line[line_addr][194] & (~hit)) | (cache_line[k][194] & (hit));
				cache_line[k][195] = (mem_line[line_addr][195] & (~hit)) | (cache_line[k][195] & (hit));
				cache_line[k][196] = (mem_line[line_addr][196] & (~hit)) | (cache_line[k][196] & (hit));
				cache_line[k][197] = (mem_line[line_addr][197] & (~hit)) | (cache_line[k][197] & (hit));
				cache_line[k][198] = (mem_line[line_addr][198] & (~hit)) | (cache_line[k][198] & (hit));
				cache_line[k][199] = (mem_line[line_addr][199] & (~hit)) | (cache_line[k][199] & (hit));
				cache_line[k][200] = (mem_line[line_addr][200] & (~hit)) | (cache_line[k][200] & (hit));
				cache_line[k][201] = (mem_line[line_addr][201] & (~hit)) | (cache_line[k][201] & (hit));
				cache_line[k][202] = (mem_line[line_addr][202] & (~hit)) | (cache_line[k][202] & (hit));
				cache_line[k][203] = (mem_line[line_addr][203] & (~hit)) | (cache_line[k][203] & (hit));
				cache_line[k][204] = (mem_line[line_addr][204] & (~hit)) | (cache_line[k][204] & (hit));
				cache_line[k][205] = (mem_line[line_addr][205] & (~hit)) | (cache_line[k][205] & (hit));
				cache_line[k][206] = (mem_line[line_addr][206] & (~hit)) | (cache_line[k][206] & (hit));
				cache_line[k][207] = (mem_line[line_addr][207] & (~hit)) | (cache_line[k][207] & (hit));
				cache_line[k][208] = (mem_line[line_addr][208] & (~hit)) | (cache_line[k][208] & (hit));
				cache_line[k][209] = (mem_line[line_addr][209] & (~hit)) | (cache_line[k][209] & (hit));
				cache_line[k][210] = (mem_line[line_addr][210] & (~hit)) | (cache_line[k][210] & (hit));
				cache_line[k][211] = (mem_line[line_addr][211] & (~hit)) | (cache_line[k][211] & (hit));
				cache_line[k][212] = (mem_line[line_addr][212] & (~hit)) | (cache_line[k][212] & (hit));
				cache_line[k][213] = (mem_line[line_addr][213] & (~hit)) | (cache_line[k][213] & (hit));
				cache_line[k][214] = (mem_line[line_addr][214] & (~hit)) | (cache_line[k][214] & (hit));
				cache_line[k][215] = (mem_line[line_addr][215] & (~hit)) | (cache_line[k][215] & (hit));
				cache_line[k][216] = (mem_line[line_addr][216] & (~hit)) | (cache_line[k][216] & (hit));
				cache_line[k][217] = (mem_line[line_addr][217] & (~hit)) | (cache_line[k][217] & (hit));
				cache_line[k][218] = (mem_line[line_addr][218] & (~hit)) | (cache_line[k][218] & (hit));
				cache_line[k][219] = (mem_line[line_addr][219] & (~hit)) | (cache_line[k][219] & (hit));
				cache_line[k][220] = (mem_line[line_addr][220] & (~hit)) | (cache_line[k][220] & (hit));
				cache_line[k][221] = (mem_line[line_addr][221] & (~hit)) | (cache_line[k][221] & (hit));
				cache_line[k][222] = (mem_line[line_addr][222] & (~hit)) | (cache_line[k][222] & (hit));
				cache_line[k][223] = (mem_line[line_addr][223] & (~hit)) | (cache_line[k][223] & (hit));
				cache_line[k][224] = (mem_line[line_addr][224] & (~hit)) | (cache_line[k][224] & (hit));
				cache_line[k][225] = (mem_line[line_addr][225] & (~hit)) | (cache_line[k][225] & (hit));
				cache_line[k][226] = (mem_line[line_addr][226] & (~hit)) | (cache_line[k][226] & (hit));
				cache_line[k][227] = (mem_line[line_addr][227] & (~hit)) | (cache_line[k][227] & (hit));
				cache_line[k][228] = (mem_line[line_addr][228] & (~hit)) | (cache_line[k][228] & (hit));
				cache_line[k][229] = (mem_line[line_addr][229] & (~hit)) | (cache_line[k][229] & (hit));
				cache_line[k][230] = (mem_line[line_addr][230] & (~hit)) | (cache_line[k][230] & (hit));
				cache_line[k][231] = (mem_line[line_addr][231] & (~hit)) | (cache_line[k][231] & (hit));
				cache_line[k][232] = (mem_line[line_addr][232] & (~hit)) | (cache_line[k][232] & (hit));
				cache_line[k][233] = (mem_line[line_addr][233] & (~hit)) | (cache_line[k][233] & (hit));
				cache_line[k][234] = (mem_line[line_addr][234] & (~hit)) | (cache_line[k][234] & (hit));
				cache_line[k][235] = (mem_line[line_addr][235] & (~hit)) | (cache_line[k][235] & (hit));
				cache_line[k][236] = (mem_line[line_addr][236] & (~hit)) | (cache_line[k][236] & (hit));
				cache_line[k][237] = (mem_line[line_addr][237] & (~hit)) | (cache_line[k][237] & (hit));
				cache_line[k][238] = (mem_line[line_addr][238] & (~hit)) | (cache_line[k][238] & (hit));
				cache_line[k][239] = (mem_line[line_addr][239] & (~hit)) | (cache_line[k][239] & (hit));
				cache_line[k][240] = (mem_line[line_addr][240] & (~hit)) | (cache_line[k][240] & (hit));
				cache_line[k][241] = (mem_line[line_addr][241] & (~hit)) | (cache_line[k][241] & (hit));
				cache_line[k][242] = (mem_line[line_addr][242] & (~hit)) | (cache_line[k][242] & (hit));
				cache_line[k][243] = (mem_line[line_addr][243] & (~hit)) | (cache_line[k][243] & (hit));
				cache_line[k][244] = (mem_line[line_addr][244] & (~hit)) | (cache_line[k][244] & (hit));
				cache_line[k][245] = (mem_line[line_addr][245] & (~hit)) | (cache_line[k][245] & (hit));
				cache_line[k][246] = (mem_line[line_addr][246] & (~hit)) | (cache_line[k][246] & (hit));
				cache_line[k][247] = (mem_line[line_addr][247] & (~hit)) | (cache_line[k][247] & (hit));
				cache_line[k][248] = (mem_line[line_addr][248] & (~hit)) | (cache_line[k][248] & (hit));
				cache_line[k][249] = (mem_line[line_addr][249] & (~hit)) | (cache_line[k][249] & (hit));
				cache_line[k][250] = (mem_line[line_addr][250] & (~hit)) | (cache_line[k][250] & (hit));
				cache_line[k][251] = (mem_line[line_addr][251] & (~hit)) | (cache_line[k][251] & (hit));
				cache_line[k][252] = (mem_line[line_addr][252] & (~hit)) | (cache_line[k][252] & (hit));
				cache_line[k][253] = (mem_line[line_addr][253] & (~hit)) | (cache_line[k][253] & (hit));
				cache_line[k][254] = (mem_line[line_addr][254] & (~hit)) | (cache_line[k][254] & (hit));
				cache_line[k][255] = (mem_line[line_addr][255] & (~hit)) | (cache_line[k][255] & (hit));
				cache_line[k][256] = (mem_line[line_addr][256] & (~hit)) | (cache_line[k][256] & (hit));
				cache_line[k][257] = (mem_line[line_addr][257] & (~hit)) | (cache_line[k][257] & (hit));
				cache_line[k][258] = (mem_line[line_addr][258] & (~hit)) | (cache_line[k][258] & (hit));
				cache_line[k][259] = (mem_line[line_addr][259] & (~hit)) | (cache_line[k][259] & (hit));
				cache_line[k][260] = (mem_line[line_addr][260] & (~hit)) | (cache_line[k][260] & (hit));
				cache_line[k][261] = (mem_line[line_addr][261] & (~hit)) | (cache_line[k][261] & (hit));
				cache_line[k][262] = (mem_line[line_addr][262] & (~hit)) | (cache_line[k][262] & (hit));
				cache_line[k][263] = (mem_line[line_addr][263] & (~hit)) | (cache_line[k][263] & (hit));
				cache_line[k][264] = (mem_line[line_addr][264] & (~hit)) | (cache_line[k][264] & (hit));
				cache_line[k][265] = (mem_line[line_addr][265] & (~hit)) | (cache_line[k][265] & (hit));
				cache_line[k][266] = (mem_line[line_addr][266] & (~hit)) | (cache_line[k][266] & (hit));
				cache_line[k][267] = (mem_line[line_addr][267] & (~hit)) | (cache_line[k][267] & (hit));
				cache_line[k][268] = (mem_line[line_addr][268] & (~hit)) | (cache_line[k][268] & (hit));
				cache_line[k][269] = (mem_line[line_addr][269] & (~hit)) | (cache_line[k][269] & (hit));
				cache_line[k][270] = (mem_line[line_addr][270] & (~hit)) | (cache_line[k][270] & (hit));
				cache_line[k][271] = (mem_line[line_addr][271] & (~hit)) | (cache_line[k][271] & (hit));
				cache_line[k][272] = (mem_line[line_addr][272] & (~hit)) | (cache_line[k][272] & (hit));
				cache_line[k][273] = (mem_line[line_addr][273] & (~hit)) | (cache_line[k][273] & (hit));
				cache_line[k][274] = (mem_line[line_addr][274] & (~hit)) | (cache_line[k][274] & (hit));
				cache_line[k][275] = (mem_line[line_addr][275] & (~hit)) | (cache_line[k][275] & (hit));
				cache_line[k][276] = (mem_line[line_addr][276] & (~hit)) | (cache_line[k][276] & (hit));
				cache_line[k][277] = (mem_line[line_addr][277] & (~hit)) | (cache_line[k][277] & (hit));
				cache_line[k][278] = (mem_line[line_addr][278] & (~hit)) | (cache_line[k][278] & (hit));
				cache_line[k][279] = (mem_line[line_addr][279] & (~hit)) | (cache_line[k][279] & (hit));
				cache_line[k][280] = (mem_line[line_addr][280] & (~hit)) | (cache_line[k][280] & (hit));
				cache_line[k][281] = (mem_line[line_addr][281] & (~hit)) | (cache_line[k][281] & (hit));
				cache_line[k][282] = (mem_line[line_addr][282] & (~hit)) | (cache_line[k][282] & (hit));
				cache_line[k][283] = (mem_line[line_addr][283] & (~hit)) | (cache_line[k][283] & (hit));
				cache_line[k][284] = (mem_line[line_addr][284] & (~hit)) | (cache_line[k][284] & (hit));
				cache_line[k][285] = (mem_line[line_addr][285] & (~hit)) | (cache_line[k][285] & (hit));
				cache_line[k][286] = (mem_line[line_addr][286] & (~hit)) | (cache_line[k][286] & (hit));
				cache_line[k][287] = (mem_line[line_addr][287] & (~hit)) | (cache_line[k][287] & (hit));
				cache_line[k][288] = (mem_line[line_addr][288] & (~hit)) | (cache_line[k][288] & (hit));
				cache_line[k][289] = (mem_line[line_addr][289] & (~hit)) | (cache_line[k][289] & (hit));
				cache_line[k][290] = (mem_line[line_addr][290] & (~hit)) | (cache_line[k][290] & (hit));
				cache_line[k][291] = (mem_line[line_addr][291] & (~hit)) | (cache_line[k][291] & (hit));
				cache_line[k][292] = (mem_line[line_addr][292] & (~hit)) | (cache_line[k][292] & (hit));
				cache_line[k][293] = (mem_line[line_addr][293] & (~hit)) | (cache_line[k][293] & (hit));
				cache_line[k][294] = (mem_line[line_addr][294] & (~hit)) | (cache_line[k][294] & (hit));
				cache_line[k][295] = (mem_line[line_addr][295] & (~hit)) | (cache_line[k][295] & (hit));
				cache_line[k][296] = (mem_line[line_addr][296] & (~hit)) | (cache_line[k][296] & (hit));
				cache_line[k][297] = (mem_line[line_addr][297] & (~hit)) | (cache_line[k][297] & (hit));
				cache_line[k][298] = (mem_line[line_addr][298] & (~hit)) | (cache_line[k][298] & (hit));
				cache_line[k][299] = (mem_line[line_addr][299] & (~hit)) | (cache_line[k][299] & (hit));
				cache_line[k][300] = (mem_line[line_addr][300] & (~hit)) | (cache_line[k][300] & (hit));
				cache_line[k][301] = (mem_line[line_addr][301] & (~hit)) | (cache_line[k][301] & (hit));
				cache_line[k][302] = (mem_line[line_addr][302] & (~hit)) | (cache_line[k][302] & (hit));
				cache_line[k][303] = (mem_line[line_addr][303] & (~hit)) | (cache_line[k][303] & (hit));
				cache_line[k][304] = (mem_line[line_addr][304] & (~hit)) | (cache_line[k][304] & (hit));
				cache_line[k][305] = (mem_line[line_addr][305] & (~hit)) | (cache_line[k][305] & (hit));
				cache_line[k][306] = (mem_line[line_addr][306] & (~hit)) | (cache_line[k][306] & (hit));
				cache_line[k][307] = (mem_line[line_addr][307] & (~hit)) | (cache_line[k][307] & (hit));
				cache_line[k][308] = (mem_line[line_addr][308] & (~hit)) | (cache_line[k][308] & (hit));
				cache_line[k][309] = (mem_line[line_addr][309] & (~hit)) | (cache_line[k][309] & (hit));
				cache_line[k][310] = (mem_line[line_addr][310] & (~hit)) | (cache_line[k][310] & (hit));
				cache_line[k][311] = (mem_line[line_addr][311] & (~hit)) | (cache_line[k][311] & (hit));
				cache_line[k][312] = (mem_line[line_addr][312] & (~hit)) | (cache_line[k][312] & (hit));
				cache_line[k][313] = (mem_line[line_addr][313] & (~hit)) | (cache_line[k][313] & (hit));
				cache_line[k][314] = (mem_line[line_addr][314] & (~hit)) | (cache_line[k][314] & (hit));
				cache_line[k][315] = (mem_line[line_addr][315] & (~hit)) | (cache_line[k][315] & (hit));
				cache_line[k][316] = (mem_line[line_addr][316] & (~hit)) | (cache_line[k][316] & (hit));
				cache_line[k][317] = (mem_line[line_addr][317] & (~hit)) | (cache_line[k][317] & (hit));
				cache_line[k][318] = (mem_line[line_addr][318] & (~hit)) | (cache_line[k][318] & (hit));
				cache_line[k][319] = (mem_line[line_addr][319] & (~hit)) | (cache_line[k][319] & (hit));
				cache_line[k][320] = (mem_line[line_addr][320] & (~hit)) | (cache_line[k][320] & (hit));
				cache_line[k][321] = (mem_line[line_addr][321] & (~hit)) | (cache_line[k][321] & (hit));
				cache_line[k][322] = (mem_line[line_addr][322] & (~hit)) | (cache_line[k][322] & (hit));
				cache_line[k][323] = (mem_line[line_addr][323] & (~hit)) | (cache_line[k][323] & (hit));
				cache_line[k][324] = (mem_line[line_addr][324] & (~hit)) | (cache_line[k][324] & (hit));
				cache_line[k][325] = (mem_line[line_addr][325] & (~hit)) | (cache_line[k][325] & (hit));
				cache_line[k][326] = (mem_line[line_addr][326] & (~hit)) | (cache_line[k][326] & (hit));
				cache_line[k][327] = (mem_line[line_addr][327] & (~hit)) | (cache_line[k][327] & (hit));
				cache_line[k][328] = (mem_line[line_addr][328] & (~hit)) | (cache_line[k][328] & (hit));
				cache_line[k][329] = (mem_line[line_addr][329] & (~hit)) | (cache_line[k][329] & (hit));
				cache_line[k][330] = (mem_line[line_addr][330] & (~hit)) | (cache_line[k][330] & (hit));
				cache_line[k][331] = (mem_line[line_addr][331] & (~hit)) | (cache_line[k][331] & (hit));
				cache_line[k][332] = (mem_line[line_addr][332] & (~hit)) | (cache_line[k][332] & (hit));
				cache_line[k][333] = (mem_line[line_addr][333] & (~hit)) | (cache_line[k][333] & (hit));
				cache_line[k][334] = (mem_line[line_addr][334] & (~hit)) | (cache_line[k][334] & (hit));
				cache_line[k][335] = (mem_line[line_addr][335] & (~hit)) | (cache_line[k][335] & (hit));
				cache_line[k][336] = (mem_line[line_addr][336] & (~hit)) | (cache_line[k][336] & (hit));
				cache_line[k][337] = (mem_line[line_addr][337] & (~hit)) | (cache_line[k][337] & (hit));
				cache_line[k][338] = (mem_line[line_addr][338] & (~hit)) | (cache_line[k][338] & (hit));
				cache_line[k][339] = (mem_line[line_addr][339] & (~hit)) | (cache_line[k][339] & (hit));
				cache_line[k][340] = (mem_line[line_addr][340] & (~hit)) | (cache_line[k][340] & (hit));
				cache_line[k][341] = (mem_line[line_addr][341] & (~hit)) | (cache_line[k][341] & (hit));
				cache_line[k][342] = (mem_line[line_addr][342] & (~hit)) | (cache_line[k][342] & (hit));
				cache_line[k][343] = (mem_line[line_addr][343] & (~hit)) | (cache_line[k][343] & (hit));
				cache_line[k][344] = (mem_line[line_addr][344] & (~hit)) | (cache_line[k][344] & (hit));
				cache_line[k][345] = (mem_line[line_addr][345] & (~hit)) | (cache_line[k][345] & (hit));
				cache_line[k][346] = (mem_line[line_addr][346] & (~hit)) | (cache_line[k][346] & (hit));
				cache_line[k][347] = (mem_line[line_addr][347] & (~hit)) | (cache_line[k][347] & (hit));
				cache_line[k][348] = (mem_line[line_addr][348] & (~hit)) | (cache_line[k][348] & (hit));
				cache_line[k][349] = (mem_line[line_addr][349] & (~hit)) | (cache_line[k][349] & (hit));
				cache_line[k][350] = (mem_line[line_addr][350] & (~hit)) | (cache_line[k][350] & (hit));
				cache_line[k][351] = (mem_line[line_addr][351] & (~hit)) | (cache_line[k][351] & (hit));
				cache_line[k][352] = (mem_line[line_addr][352] & (~hit)) | (cache_line[k][352] & (hit));
				cache_line[k][353] = (mem_line[line_addr][353] & (~hit)) | (cache_line[k][353] & (hit));
				cache_line[k][354] = (mem_line[line_addr][354] & (~hit)) | (cache_line[k][354] & (hit));
				cache_line[k][355] = (mem_line[line_addr][355] & (~hit)) | (cache_line[k][355] & (hit));
				cache_line[k][356] = (mem_line[line_addr][356] & (~hit)) | (cache_line[k][356] & (hit));
				cache_line[k][357] = (mem_line[line_addr][357] & (~hit)) | (cache_line[k][357] & (hit));
				cache_line[k][358] = (mem_line[line_addr][358] & (~hit)) | (cache_line[k][358] & (hit));
				cache_line[k][359] = (mem_line[line_addr][359] & (~hit)) | (cache_line[k][359] & (hit));
				cache_line[k][360] = (mem_line[line_addr][360] & (~hit)) | (cache_line[k][360] & (hit));
				cache_line[k][361] = (mem_line[line_addr][361] & (~hit)) | (cache_line[k][361] & (hit));
				cache_line[k][362] = (mem_line[line_addr][362] & (~hit)) | (cache_line[k][362] & (hit));
				cache_line[k][363] = (mem_line[line_addr][363] & (~hit)) | (cache_line[k][363] & (hit));
				cache_line[k][364] = (mem_line[line_addr][364] & (~hit)) | (cache_line[k][364] & (hit));
				cache_line[k][365] = (mem_line[line_addr][365] & (~hit)) | (cache_line[k][365] & (hit));
				cache_line[k][366] = (mem_line[line_addr][366] & (~hit)) | (cache_line[k][366] & (hit));
				cache_line[k][367] = (mem_line[line_addr][367] & (~hit)) | (cache_line[k][367] & (hit));
				cache_line[k][368] = (mem_line[line_addr][368] & (~hit)) | (cache_line[k][368] & (hit));
				cache_line[k][369] = (mem_line[line_addr][369] & (~hit)) | (cache_line[k][369] & (hit));
				cache_line[k][370] = (mem_line[line_addr][370] & (~hit)) | (cache_line[k][370] & (hit));
				cache_line[k][371] = (mem_line[line_addr][371] & (~hit)) | (cache_line[k][371] & (hit));
				cache_line[k][372] = (mem_line[line_addr][372] & (~hit)) | (cache_line[k][372] & (hit));
				cache_line[k][373] = (mem_line[line_addr][373] & (~hit)) | (cache_line[k][373] & (hit));
				cache_line[k][374] = (mem_line[line_addr][374] & (~hit)) | (cache_line[k][374] & (hit));
				cache_line[k][375] = (mem_line[line_addr][375] & (~hit)) | (cache_line[k][375] & (hit));
				cache_line[k][376] = (mem_line[line_addr][376] & (~hit)) | (cache_line[k][376] & (hit));
				cache_line[k][377] = (mem_line[line_addr][377] & (~hit)) | (cache_line[k][377] & (hit));
				cache_line[k][378] = (mem_line[line_addr][378] & (~hit)) | (cache_line[k][378] & (hit));
				cache_line[k][379] = (mem_line[line_addr][379] & (~hit)) | (cache_line[k][379] & (hit));
				cache_line[k][380] = (mem_line[line_addr][380] & (~hit)) | (cache_line[k][380] & (hit));
				cache_line[k][381] = (mem_line[line_addr][381] & (~hit)) | (cache_line[k][381] & (hit));
				cache_line[k][382] = (mem_line[line_addr][382] & (~hit)) | (cache_line[k][382] & (hit));
				cache_line[k][383] = (mem_line[line_addr][383] & (~hit)) | (cache_line[k][383] & (hit));
				cache_line[k][384] = (mem_line[line_addr][384] & (~hit)) | (cache_line[k][384] & (hit));
				cache_line[k][385] = (mem_line[line_addr][385] & (~hit)) | (cache_line[k][385] & (hit));
				cache_line[k][386] = (mem_line[line_addr][386] & (~hit)) | (cache_line[k][386] & (hit));
				cache_line[k][387] = (mem_line[line_addr][387] & (~hit)) | (cache_line[k][387] & (hit));
				cache_line[k][388] = (mem_line[line_addr][388] & (~hit)) | (cache_line[k][388] & (hit));
				cache_line[k][389] = (mem_line[line_addr][389] & (~hit)) | (cache_line[k][389] & (hit));
				cache_line[k][390] = (mem_line[line_addr][390] & (~hit)) | (cache_line[k][390] & (hit));
				cache_line[k][391] = (mem_line[line_addr][391] & (~hit)) | (cache_line[k][391] & (hit));
				cache_line[k][392] = (mem_line[line_addr][392] & (~hit)) | (cache_line[k][392] & (hit));
				cache_line[k][393] = (mem_line[line_addr][393] & (~hit)) | (cache_line[k][393] & (hit));
				cache_line[k][394] = (mem_line[line_addr][394] & (~hit)) | (cache_line[k][394] & (hit));
				cache_line[k][395] = (mem_line[line_addr][395] & (~hit)) | (cache_line[k][395] & (hit));
				cache_line[k][396] = (mem_line[line_addr][396] & (~hit)) | (cache_line[k][396] & (hit));
				cache_line[k][397] = (mem_line[line_addr][397] & (~hit)) | (cache_line[k][397] & (hit));
				cache_line[k][398] = (mem_line[line_addr][398] & (~hit)) | (cache_line[k][398] & (hit));
				cache_line[k][399] = (mem_line[line_addr][399] & (~hit)) | (cache_line[k][399] & (hit));
				cache_line[k][400] = (mem_line[line_addr][400] & (~hit)) | (cache_line[k][400] & (hit));
				cache_line[k][401] = (mem_line[line_addr][401] & (~hit)) | (cache_line[k][401] & (hit));
				cache_line[k][402] = (mem_line[line_addr][402] & (~hit)) | (cache_line[k][402] & (hit));
				cache_line[k][403] = (mem_line[line_addr][403] & (~hit)) | (cache_line[k][403] & (hit));
				cache_line[k][404] = (mem_line[line_addr][404] & (~hit)) | (cache_line[k][404] & (hit));
				cache_line[k][405] = (mem_line[line_addr][405] & (~hit)) | (cache_line[k][405] & (hit));
				cache_line[k][406] = (mem_line[line_addr][406] & (~hit)) | (cache_line[k][406] & (hit));
				cache_line[k][407] = (mem_line[line_addr][407] & (~hit)) | (cache_line[k][407] & (hit));
				cache_line[k][408] = (mem_line[line_addr][408] & (~hit)) | (cache_line[k][408] & (hit));
				cache_line[k][409] = (mem_line[line_addr][409] & (~hit)) | (cache_line[k][409] & (hit));
				cache_line[k][410] = (mem_line[line_addr][410] & (~hit)) | (cache_line[k][410] & (hit));
				cache_line[k][411] = (mem_line[line_addr][411] & (~hit)) | (cache_line[k][411] & (hit));
				cache_line[k][412] = (mem_line[line_addr][412] & (~hit)) | (cache_line[k][412] & (hit));
				cache_line[k][413] = (mem_line[line_addr][413] & (~hit)) | (cache_line[k][413] & (hit));
				cache_line[k][414] = (mem_line[line_addr][414] & (~hit)) | (cache_line[k][414] & (hit));
				cache_line[k][415] = (mem_line[line_addr][415] & (~hit)) | (cache_line[k][415] & (hit));
				cache_line[k][416] = (mem_line[line_addr][416] & (~hit)) | (cache_line[k][416] & (hit));
				cache_line[k][417] = (mem_line[line_addr][417] & (~hit)) | (cache_line[k][417] & (hit));
				cache_line[k][418] = (mem_line[line_addr][418] & (~hit)) | (cache_line[k][418] & (hit));
				cache_line[k][419] = (mem_line[line_addr][419] & (~hit)) | (cache_line[k][419] & (hit));
				cache_line[k][420] = (mem_line[line_addr][420] & (~hit)) | (cache_line[k][420] & (hit));
				cache_line[k][421] = (mem_line[line_addr][421] & (~hit)) | (cache_line[k][421] & (hit));
				cache_line[k][422] = (mem_line[line_addr][422] & (~hit)) | (cache_line[k][422] & (hit));
				cache_line[k][423] = (mem_line[line_addr][423] & (~hit)) | (cache_line[k][423] & (hit));
				cache_line[k][424] = (mem_line[line_addr][424] & (~hit)) | (cache_line[k][424] & (hit));
				cache_line[k][425] = (mem_line[line_addr][425] & (~hit)) | (cache_line[k][425] & (hit));
				cache_line[k][426] = (mem_line[line_addr][426] & (~hit)) | (cache_line[k][426] & (hit));
				cache_line[k][427] = (mem_line[line_addr][427] & (~hit)) | (cache_line[k][427] & (hit));
				cache_line[k][428] = (mem_line[line_addr][428] & (~hit)) | (cache_line[k][428] & (hit));
				cache_line[k][429] = (mem_line[line_addr][429] & (~hit)) | (cache_line[k][429] & (hit));
				cache_line[k][430] = (mem_line[line_addr][430] & (~hit)) | (cache_line[k][430] & (hit));
				cache_line[k][431] = (mem_line[line_addr][431] & (~hit)) | (cache_line[k][431] & (hit));
				cache_line[k][432] = (mem_line[line_addr][432] & (~hit)) | (cache_line[k][432] & (hit));
				cache_line[k][433] = (mem_line[line_addr][433] & (~hit)) | (cache_line[k][433] & (hit));
				cache_line[k][434] = (mem_line[line_addr][434] & (~hit)) | (cache_line[k][434] & (hit));
				cache_line[k][435] = (mem_line[line_addr][435] & (~hit)) | (cache_line[k][435] & (hit));
				cache_line[k][436] = (mem_line[line_addr][436] & (~hit)) | (cache_line[k][436] & (hit));
				cache_line[k][437] = (mem_line[line_addr][437] & (~hit)) | (cache_line[k][437] & (hit));
				cache_line[k][438] = (mem_line[line_addr][438] & (~hit)) | (cache_line[k][438] & (hit));
				cache_line[k][439] = (mem_line[line_addr][439] & (~hit)) | (cache_line[k][439] & (hit));
				cache_line[k][440] = (mem_line[line_addr][440] & (~hit)) | (cache_line[k][440] & (hit));
				cache_line[k][441] = (mem_line[line_addr][441] & (~hit)) | (cache_line[k][441] & (hit));
				cache_line[k][442] = (mem_line[line_addr][442] & (~hit)) | (cache_line[k][442] & (hit));
				cache_line[k][443] = (mem_line[line_addr][443] & (~hit)) | (cache_line[k][443] & (hit));
				cache_line[k][444] = (mem_line[line_addr][444] & (~hit)) | (cache_line[k][444] & (hit));
				cache_line[k][445] = (mem_line[line_addr][445] & (~hit)) | (cache_line[k][445] & (hit));
				cache_line[k][446] = (mem_line[line_addr][446] & (~hit)) | (cache_line[k][446] & (hit));
				cache_line[k][447] = (mem_line[line_addr][447] & (~hit)) | (cache_line[k][447] & (hit));
				cache_line[k][448] = (mem_line[line_addr][448] & (~hit)) | (cache_line[k][448] & (hit));
				cache_line[k][449] = (mem_line[line_addr][449] & (~hit)) | (cache_line[k][449] & (hit));
				cache_line[k][450] = (mem_line[line_addr][450] & (~hit)) | (cache_line[k][450] & (hit));
				cache_line[k][451] = (mem_line[line_addr][451] & (~hit)) | (cache_line[k][451] & (hit));
				cache_line[k][452] = (mem_line[line_addr][452] & (~hit)) | (cache_line[k][452] & (hit));
				cache_line[k][453] = (mem_line[line_addr][453] & (~hit)) | (cache_line[k][453] & (hit));
				cache_line[k][454] = (mem_line[line_addr][454] & (~hit)) | (cache_line[k][454] & (hit));
				cache_line[k][455] = (mem_line[line_addr][455] & (~hit)) | (cache_line[k][455] & (hit));
				cache_line[k][456] = (mem_line[line_addr][456] & (~hit)) | (cache_line[k][456] & (hit));
				cache_line[k][457] = (mem_line[line_addr][457] & (~hit)) | (cache_line[k][457] & (hit));
				cache_line[k][458] = (mem_line[line_addr][458] & (~hit)) | (cache_line[k][458] & (hit));
				cache_line[k][459] = (mem_line[line_addr][459] & (~hit)) | (cache_line[k][459] & (hit));
				cache_line[k][460] = (mem_line[line_addr][460] & (~hit)) | (cache_line[k][460] & (hit));
				cache_line[k][461] = (mem_line[line_addr][461] & (~hit)) | (cache_line[k][461] & (hit));
				cache_line[k][462] = (mem_line[line_addr][462] & (~hit)) | (cache_line[k][462] & (hit));
				cache_line[k][463] = (mem_line[line_addr][463] & (~hit)) | (cache_line[k][463] & (hit));
				cache_line[k][464] = (mem_line[line_addr][464] & (~hit)) | (cache_line[k][464] & (hit));
				cache_line[k][465] = (mem_line[line_addr][465] & (~hit)) | (cache_line[k][465] & (hit));
				cache_line[k][466] = (mem_line[line_addr][466] & (~hit)) | (cache_line[k][466] & (hit));
				cache_line[k][467] = (mem_line[line_addr][467] & (~hit)) | (cache_line[k][467] & (hit));
				cache_line[k][468] = (mem_line[line_addr][468] & (~hit)) | (cache_line[k][468] & (hit));
				cache_line[k][469] = (mem_line[line_addr][469] & (~hit)) | (cache_line[k][469] & (hit));
				cache_line[k][470] = (mem_line[line_addr][470] & (~hit)) | (cache_line[k][470] & (hit));
				cache_line[k][471] = (mem_line[line_addr][471] & (~hit)) | (cache_line[k][471] & (hit));
				cache_line[k][472] = (mem_line[line_addr][472] & (~hit)) | (cache_line[k][472] & (hit));
				cache_line[k][473] = (mem_line[line_addr][473] & (~hit)) | (cache_line[k][473] & (hit));
				cache_line[k][474] = (mem_line[line_addr][474] & (~hit)) | (cache_line[k][474] & (hit));
				cache_line[k][475] = (mem_line[line_addr][475] & (~hit)) | (cache_line[k][475] & (hit));
				cache_line[k][476] = (mem_line[line_addr][476] & (~hit)) | (cache_line[k][476] & (hit));
				cache_line[k][477] = (mem_line[line_addr][477] & (~hit)) | (cache_line[k][477] & (hit));
				cache_line[k][478] = (mem_line[line_addr][478] & (~hit)) | (cache_line[k][478] & (hit));
				cache_line[k][479] = (mem_line[line_addr][479] & (~hit)) | (cache_line[k][479] & (hit));
				cache_line[k][480] = (mem_line[line_addr][480] & (~hit)) | (cache_line[k][480] & (hit));
				cache_line[k][481] = (mem_line[line_addr][481] & (~hit)) | (cache_line[k][481] & (hit));
				cache_line[k][482] = (mem_line[line_addr][482] & (~hit)) | (cache_line[k][482] & (hit));
				cache_line[k][483] = (mem_line[line_addr][483] & (~hit)) | (cache_line[k][483] & (hit));
				cache_line[k][484] = (mem_line[line_addr][484] & (~hit)) | (cache_line[k][484] & (hit));
				cache_line[k][485] = (mem_line[line_addr][485] & (~hit)) | (cache_line[k][485] & (hit));
				cache_line[k][486] = (mem_line[line_addr][486] & (~hit)) | (cache_line[k][486] & (hit));
				cache_line[k][487] = (mem_line[line_addr][487] & (~hit)) | (cache_line[k][487] & (hit));
				cache_line[k][488] = (mem_line[line_addr][488] & (~hit)) | (cache_line[k][488] & (hit));
				cache_line[k][489] = (mem_line[line_addr][489] & (~hit)) | (cache_line[k][489] & (hit));
				cache_line[k][490] = (mem_line[line_addr][490] & (~hit)) | (cache_line[k][490] & (hit));
				cache_line[k][491] = (mem_line[line_addr][491] & (~hit)) | (cache_line[k][491] & (hit));
				cache_line[k][492] = (mem_line[line_addr][492] & (~hit)) | (cache_line[k][492] & (hit));
				cache_line[k][493] = (mem_line[line_addr][493] & (~hit)) | (cache_line[k][493] & (hit));
				cache_line[k][494] = (mem_line[line_addr][494] & (~hit)) | (cache_line[k][494] & (hit));
				cache_line[k][495] = (mem_line[line_addr][495] & (~hit)) | (cache_line[k][495] & (hit));
				cache_line[k][496] = (mem_line[line_addr][496] & (~hit)) | (cache_line[k][496] & (hit));
				cache_line[k][497] = (mem_line[line_addr][497] & (~hit)) | (cache_line[k][497] & (hit));
				cache_line[k][498] = (mem_line[line_addr][498] & (~hit)) | (cache_line[k][498] & (hit));
				cache_line[k][499] = (mem_line[line_addr][499] & (~hit)) | (cache_line[k][499] & (hit));
				cache_line[k][500] = (mem_line[line_addr][500] & (~hit)) | (cache_line[k][500] & (hit));
				cache_line[k][501] = (mem_line[line_addr][501] & (~hit)) | (cache_line[k][501] & (hit));
				cache_line[k][502] = (mem_line[line_addr][502] & (~hit)) | (cache_line[k][502] & (hit));
				cache_line[k][503] = (mem_line[line_addr][503] & (~hit)) | (cache_line[k][503] & (hit));
				cache_line[k][504] = (mem_line[line_addr][504] & (~hit)) | (cache_line[k][504] & (hit));
				cache_line[k][505] = (mem_line[line_addr][505] & (~hit)) | (cache_line[k][505] & (hit));
				cache_line[k][506] = (mem_line[line_addr][506] & (~hit)) | (cache_line[k][506] & (hit));
				cache_line[k][507] = (mem_line[line_addr][507] & (~hit)) | (cache_line[k][507] & (hit));
				cache_line[k][508] = (mem_line[line_addr][508] & (~hit)) | (cache_line[k][508] & (hit));
				cache_line[k][509] = (mem_line[line_addr][509] & (~hit)) | (cache_line[k][509] & (hit));
				cache_line[k][510] = (mem_line[line_addr][510] & (~hit)) | (cache_line[k][510] & (hit));
				cache_line[k][511] = (mem_line[line_addr][511] & (~hit)) | (cache_line[k][511] & (hit));
				cache_line[k][512] = (mem_line[line_addr][512] & (~hit)) | (cache_line[k][512] & (hit));
				cache_line[k][513] = (mem_line[line_addr][513] & (~hit)) | (cache_line[k][513] & (hit));
				cache_line[k][514] = (mem_line[line_addr][514] & (~hit)) | (cache_line[k][514] & (hit));
				cache_line[k][515] = (mem_line[line_addr][515] & (~hit)) | (cache_line[k][515] & (hit));
				cache_line[k][516] = (mem_line[line_addr][516] & (~hit)) | (cache_line[k][516] & (hit));
				cache_line[k][517] = (mem_line[line_addr][517] & (~hit)) | (cache_line[k][517] & (hit));
				cache_line[k][518] = (mem_line[line_addr][518] & (~hit)) | (cache_line[k][518] & (hit));
				cache_line[k][519] = (mem_line[line_addr][519] & (~hit)) | (cache_line[k][519] & (hit));
				cache_line[k][520] = (mem_line[line_addr][520] & (~hit)) | (cache_line[k][520] & (hit));
				cache_line[k][521] = (mem_line[line_addr][521] & (~hit)) | (cache_line[k][521] & (hit));
				cache_line[k][522] = (mem_line[line_addr][522] & (~hit)) | (cache_line[k][522] & (hit));
				cache_line[k][523] = (mem_line[line_addr][523] & (~hit)) | (cache_line[k][523] & (hit));
				cache_line[k][524] = (mem_line[line_addr][524] & (~hit)) | (cache_line[k][524] & (hit));
				cache_line[k][525] = (mem_line[line_addr][525] & (~hit)) | (cache_line[k][525] & (hit));
				cache_line[k][526] = (mem_line[line_addr][526] & (~hit)) | (cache_line[k][526] & (hit));
				cache_line[k][527] = (mem_line[line_addr][527] & (~hit)) | (cache_line[k][527] & (hit));
				cache_line[k][528] = (mem_line[line_addr][528] & (~hit)) | (cache_line[k][528] & (hit));
				cache_line[k][529] = (mem_line[line_addr][529] & (~hit)) | (cache_line[k][529] & (hit));
				cache_line[k][530] = (mem_line[line_addr][530] & (~hit)) | (cache_line[k][530] & (hit));
				cache_line[k][531] = (mem_line[line_addr][531] & (~hit)) | (cache_line[k][531] & (hit));
				cache_line[k][532] = (mem_line[line_addr][532] & (~hit)) | (cache_line[k][532] & (hit));
				cache_line[k][533] = (mem_line[line_addr][533] & (~hit)) | (cache_line[k][533] & (hit));
				cache_line[k][534] = (mem_line[line_addr][534] & (~hit)) | (cache_line[k][534] & (hit));
				cache_line[k][535] = (mem_line[line_addr][535] & (~hit)) | (cache_line[k][535] & (hit));
				cache_line[k][536] = (mem_line[line_addr][536] & (~hit)) | (cache_line[k][536] & (hit));
				cache_line[k][537] = (mem_line[line_addr][537] & (~hit)) | (cache_line[k][537] & (hit));
				cache_line[k][538] = (mem_line[line_addr][538] & (~hit)) | (cache_line[k][538] & (hit));
				cache_line[k][539] = (mem_line[line_addr][539] & (~hit)) | (cache_line[k][539] & (hit));
				cache_line[k][540] = (mem_line[line_addr][540] & (~hit)) | (cache_line[k][540] & (hit));
				cache_line[k][541] = (mem_line[line_addr][541] & (~hit)) | (cache_line[k][541] & (hit));
				cache_line[k][542] = (mem_line[line_addr][542] & (~hit)) | (cache_line[k][542] & (hit));
				cache_line[k][543] = (mem_line[line_addr][543] & (~hit)) | (cache_line[k][543] & (hit));
				cache_line[k][544] = (mem_line[line_addr][544] & (~hit)) | (cache_line[k][544] & (hit));
				cache_line[k][545] = (mem_line[line_addr][545] & (~hit)) | (cache_line[k][545] & (hit));
				cache_line[k][546] = (mem_line[line_addr][546] & (~hit)) | (cache_line[k][546] & (hit));
				cache_line[k][547] = (mem_line[line_addr][547] & (~hit)) | (cache_line[k][547] & (hit));
				cache_line[k][548] = (mem_line[line_addr][548] & (~hit)) | (cache_line[k][548] & (hit));
				cache_line[k][549] = (mem_line[line_addr][549] & (~hit)) | (cache_line[k][549] & (hit));
				cache_line[k][550] = (mem_line[line_addr][550] & (~hit)) | (cache_line[k][550] & (hit));
				cache_line[k][551] = (mem_line[line_addr][551] & (~hit)) | (cache_line[k][551] & (hit));
				cache_line[k][552] = (mem_line[line_addr][552] & (~hit)) | (cache_line[k][552] & (hit));
				cache_line[k][553] = (mem_line[line_addr][553] & (~hit)) | (cache_line[k][553] & (hit));
				cache_line[k][554] = (mem_line[line_addr][554] & (~hit)) | (cache_line[k][554] & (hit));
				cache_line[k][555] = (mem_line[line_addr][555] & (~hit)) | (cache_line[k][555] & (hit));
				cache_line[k][556] = (mem_line[line_addr][556] & (~hit)) | (cache_line[k][556] & (hit));
				cache_line[k][557] = (mem_line[line_addr][557] & (~hit)) | (cache_line[k][557] & (hit));
				cache_line[k][558] = (mem_line[line_addr][558] & (~hit)) | (cache_line[k][558] & (hit));
				cache_line[k][559] = (mem_line[line_addr][559] & (~hit)) | (cache_line[k][559] & (hit));
				cache_line[k][560] = (mem_line[line_addr][560] & (~hit)) | (cache_line[k][560] & (hit));
				cache_line[k][561] = (mem_line[line_addr][561] & (~hit)) | (cache_line[k][561] & (hit));
				cache_line[k][562] = (mem_line[line_addr][562] & (~hit)) | (cache_line[k][562] & (hit));
				cache_line[k][563] = (mem_line[line_addr][563] & (~hit)) | (cache_line[k][563] & (hit));
				cache_line[k][564] = (mem_line[line_addr][564] & (~hit)) | (cache_line[k][564] & (hit));
				cache_line[k][565] = (mem_line[line_addr][565] & (~hit)) | (cache_line[k][565] & (hit));
				cache_line[k][566] = (mem_line[line_addr][566] & (~hit)) | (cache_line[k][566] & (hit));
				cache_line[k][567] = (mem_line[line_addr][567] & (~hit)) | (cache_line[k][567] & (hit));
				cache_line[k][568] = (mem_line[line_addr][568] & (~hit)) | (cache_line[k][568] & (hit));
				cache_line[k][569] = (mem_line[line_addr][569] & (~hit)) | (cache_line[k][569] & (hit));
				cache_line[k][570] = (mem_line[line_addr][570] & (~hit)) | (cache_line[k][570] & (hit));
				cache_line[k][571] = (mem_line[line_addr][571] & (~hit)) | (cache_line[k][571] & (hit));
				cache_line[k][572] = (mem_line[line_addr][572] & (~hit)) | (cache_line[k][572] & (hit));
				cache_line[k][573] = (mem_line[line_addr][573] & (~hit)) | (cache_line[k][573] & (hit));
				cache_line[k][574] = (mem_line[line_addr][574] & (~hit)) | (cache_line[k][574] & (hit));
				cache_line[k][575] = (mem_line[line_addr][575] & (~hit)) | (cache_line[k][575] & (hit));
				cache_line[k][576] = (mem_line[line_addr][576] & (~hit)) | (cache_line[k][576] & (hit));
				cache_line[k][577] = (mem_line[line_addr][577] & (~hit)) | (cache_line[k][577] & (hit));
				cache_line[k][578] = (mem_line[line_addr][578] & (~hit)) | (cache_line[k][578] & (hit));
				cache_line[k][579] = (mem_line[line_addr][579] & (~hit)) | (cache_line[k][579] & (hit));
				cache_line[k][580] = (mem_line[line_addr][580] & (~hit)) | (cache_line[k][580] & (hit));
				cache_line[k][581] = (mem_line[line_addr][581] & (~hit)) | (cache_line[k][581] & (hit));
				cache_line[k][582] = (mem_line[line_addr][582] & (~hit)) | (cache_line[k][582] & (hit));
				cache_line[k][583] = (mem_line[line_addr][583] & (~hit)) | (cache_line[k][583] & (hit));
				cache_line[k][584] = (mem_line[line_addr][584] & (~hit)) | (cache_line[k][584] & (hit));
				cache_line[k][585] = (mem_line[line_addr][585] & (~hit)) | (cache_line[k][585] & (hit));
				cache_line[k][586] = (mem_line[line_addr][586] & (~hit)) | (cache_line[k][586] & (hit));
				cache_line[k][587] = (mem_line[line_addr][587] & (~hit)) | (cache_line[k][587] & (hit));
				cache_line[k][588] = (mem_line[line_addr][588] & (~hit)) | (cache_line[k][588] & (hit));
				cache_line[k][589] = (mem_line[line_addr][589] & (~hit)) | (cache_line[k][589] & (hit));
				cache_line[k][590] = (mem_line[line_addr][590] & (~hit)) | (cache_line[k][590] & (hit));
				cache_line[k][591] = (mem_line[line_addr][591] & (~hit)) | (cache_line[k][591] & (hit));
				cache_line[k][592] = (mem_line[line_addr][592] & (~hit)) | (cache_line[k][592] & (hit));
				cache_line[k][593] = (mem_line[line_addr][593] & (~hit)) | (cache_line[k][593] & (hit));
				cache_line[k][594] = (mem_line[line_addr][594] & (~hit)) | (cache_line[k][594] & (hit));
				cache_line[k][595] = (mem_line[line_addr][595] & (~hit)) | (cache_line[k][595] & (hit));
				cache_line[k][596] = (mem_line[line_addr][596] & (~hit)) | (cache_line[k][596] & (hit));
				cache_line[k][597] = (mem_line[line_addr][597] & (~hit)) | (cache_line[k][597] & (hit));
				cache_line[k][598] = (mem_line[line_addr][598] & (~hit)) | (cache_line[k][598] & (hit));
				cache_line[k][599] = (mem_line[line_addr][599] & (~hit)) | (cache_line[k][599] & (hit));
				cache_line[k][600] = (mem_line[line_addr][600] & (~hit)) | (cache_line[k][600] & (hit));
				cache_line[k][601] = (mem_line[line_addr][601] & (~hit)) | (cache_line[k][601] & (hit));
				cache_line[k][602] = (mem_line[line_addr][602] & (~hit)) | (cache_line[k][602] & (hit));
				cache_line[k][603] = (mem_line[line_addr][603] & (~hit)) | (cache_line[k][603] & (hit));
				cache_line[k][604] = (mem_line[line_addr][604] & (~hit)) | (cache_line[k][604] & (hit));
				cache_line[k][605] = (mem_line[line_addr][605] & (~hit)) | (cache_line[k][605] & (hit));
				cache_line[k][606] = (mem_line[line_addr][606] & (~hit)) | (cache_line[k][606] & (hit));
				cache_line[k][607] = (mem_line[line_addr][607] & (~hit)) | (cache_line[k][607] & (hit));
				cache_line[k][608] = (mem_line[line_addr][608] & (~hit)) | (cache_line[k][608] & (hit));
				cache_line[k][609] = (mem_line[line_addr][609] & (~hit)) | (cache_line[k][609] & (hit));
				cache_line[k][610] = (mem_line[line_addr][610] & (~hit)) | (cache_line[k][610] & (hit));
				cache_line[k][611] = (mem_line[line_addr][611] & (~hit)) | (cache_line[k][611] & (hit));
				cache_line[k][612] = (mem_line[line_addr][612] & (~hit)) | (cache_line[k][612] & (hit));
				cache_line[k][613] = (mem_line[line_addr][613] & (~hit)) | (cache_line[k][613] & (hit));
				cache_line[k][614] = (mem_line[line_addr][614] & (~hit)) | (cache_line[k][614] & (hit));
				cache_line[k][615] = (mem_line[line_addr][615] & (~hit)) | (cache_line[k][615] & (hit));
				cache_line[k][616] = (mem_line[line_addr][616] & (~hit)) | (cache_line[k][616] & (hit));
				cache_line[k][617] = (mem_line[line_addr][617] & (~hit)) | (cache_line[k][617] & (hit));
				cache_line[k][618] = (mem_line[line_addr][618] & (~hit)) | (cache_line[k][618] & (hit));
				cache_line[k][619] = (mem_line[line_addr][619] & (~hit)) | (cache_line[k][619] & (hit));
				cache_line[k][620] = (mem_line[line_addr][620] & (~hit)) | (cache_line[k][620] & (hit));
				cache_line[k][621] = (mem_line[line_addr][621] & (~hit)) | (cache_line[k][621] & (hit));
				cache_line[k][622] = (mem_line[line_addr][622] & (~hit)) | (cache_line[k][622] & (hit));
				cache_line[k][623] = (mem_line[line_addr][623] & (~hit)) | (cache_line[k][623] & (hit));
				cache_line[k][624] = (mem_line[line_addr][624] & (~hit)) | (cache_line[k][624] & (hit));
				cache_line[k][625] = (mem_line[line_addr][625] & (~hit)) | (cache_line[k][625] & (hit));
				cache_line[k][626] = (mem_line[line_addr][626] & (~hit)) | (cache_line[k][626] & (hit));
				cache_line[k][627] = (mem_line[line_addr][627] & (~hit)) | (cache_line[k][627] & (hit));
				cache_line[k][628] = (mem_line[line_addr][628] & (~hit)) | (cache_line[k][628] & (hit));
				cache_line[k][629] = (mem_line[line_addr][629] & (~hit)) | (cache_line[k][629] & (hit));
				cache_line[k][630] = (mem_line[line_addr][630] & (~hit)) | (cache_line[k][630] & (hit));
				cache_line[k][631] = (mem_line[line_addr][631] & (~hit)) | (cache_line[k][631] & (hit));
				cache_line[k][632] = (mem_line[line_addr][632] & (~hit)) | (cache_line[k][632] & (hit));
				cache_line[k][633] = (mem_line[line_addr][633] & (~hit)) | (cache_line[k][633] & (hit));
				cache_line[k][634] = (mem_line[line_addr][634] & (~hit)) | (cache_line[k][634] & (hit));
				cache_line[k][635] = (mem_line[line_addr][635] & (~hit)) | (cache_line[k][635] & (hit));
				cache_line[k][636] = (mem_line[line_addr][636] & (~hit)) | (cache_line[k][636] & (hit));
				cache_line[k][637] = (mem_line[line_addr][637] & (~hit)) | (cache_line[k][637] & (hit));
				cache_line[k][638] = (mem_line[line_addr][638] & (~hit)) | (cache_line[k][638] & (hit));
				cache_line[k][639] = (mem_line[line_addr][639] & (~hit)) | (cache_line[k][639] & (hit));
				cache_line[k][640] = (mem_line[line_addr][640] & (~hit)) | (cache_line[k][640] & (hit));
				cache_line[k][641] = (mem_line[line_addr][641] & (~hit)) | (cache_line[k][641] & (hit));
				cache_line[k][642] = (mem_line[line_addr][642] & (~hit)) | (cache_line[k][642] & (hit));
				cache_line[k][643] = (mem_line[line_addr][643] & (~hit)) | (cache_line[k][643] & (hit));
				cache_line[k][644] = (mem_line[line_addr][644] & (~hit)) | (cache_line[k][644] & (hit));
				cache_line[k][645] = (mem_line[line_addr][645] & (~hit)) | (cache_line[k][645] & (hit));
				cache_line[k][646] = (mem_line[line_addr][646] & (~hit)) | (cache_line[k][646] & (hit));
				cache_line[k][647] = (mem_line[line_addr][647] & (~hit)) | (cache_line[k][647] & (hit));
				cache_line[k][648] = (mem_line[line_addr][648] & (~hit)) | (cache_line[k][648] & (hit));
				cache_line[k][649] = (mem_line[line_addr][649] & (~hit)) | (cache_line[k][649] & (hit));
				cache_line[k][650] = (mem_line[line_addr][650] & (~hit)) | (cache_line[k][650] & (hit));
				cache_line[k][651] = (mem_line[line_addr][651] & (~hit)) | (cache_line[k][651] & (hit));
				cache_line[k][652] = (mem_line[line_addr][652] & (~hit)) | (cache_line[k][652] & (hit));
				cache_line[k][653] = (mem_line[line_addr][653] & (~hit)) | (cache_line[k][653] & (hit));
				cache_line[k][654] = (mem_line[line_addr][654] & (~hit)) | (cache_line[k][654] & (hit));
				cache_line[k][655] = (mem_line[line_addr][655] & (~hit)) | (cache_line[k][655] & (hit));
				cache_line[k][656] = (mem_line[line_addr][656] & (~hit)) | (cache_line[k][656] & (hit));
				cache_line[k][657] = (mem_line[line_addr][657] & (~hit)) | (cache_line[k][657] & (hit));
				cache_line[k][658] = (mem_line[line_addr][658] & (~hit)) | (cache_line[k][658] & (hit));
				cache_line[k][659] = (mem_line[line_addr][659] & (~hit)) | (cache_line[k][659] & (hit));
				cache_line[k][660] = (mem_line[line_addr][660] & (~hit)) | (cache_line[k][660] & (hit));
				cache_line[k][661] = (mem_line[line_addr][661] & (~hit)) | (cache_line[k][661] & (hit));
				cache_line[k][662] = (mem_line[line_addr][662] & (~hit)) | (cache_line[k][662] & (hit));
				cache_line[k][663] = (mem_line[line_addr][663] & (~hit)) | (cache_line[k][663] & (hit));
				cache_line[k][664] = (mem_line[line_addr][664] & (~hit)) | (cache_line[k][664] & (hit));
				cache_line[k][665] = (mem_line[line_addr][665] & (~hit)) | (cache_line[k][665] & (hit));
				cache_line[k][666] = (mem_line[line_addr][666] & (~hit)) | (cache_line[k][666] & (hit));
				cache_line[k][667] = (mem_line[line_addr][667] & (~hit)) | (cache_line[k][667] & (hit));
				cache_line[k][668] = (mem_line[line_addr][668] & (~hit)) | (cache_line[k][668] & (hit));
				cache_line[k][669] = (mem_line[line_addr][669] & (~hit)) | (cache_line[k][669] & (hit));
				cache_line[k][670] = (mem_line[line_addr][670] & (~hit)) | (cache_line[k][670] & (hit));
				cache_line[k][671] = (mem_line[line_addr][671] & (~hit)) | (cache_line[k][671] & (hit));
				cache_line[k][672] = (mem_line[line_addr][672] & (~hit)) | (cache_line[k][672] & (hit));
				cache_line[k][673] = (mem_line[line_addr][673] & (~hit)) | (cache_line[k][673] & (hit));
				cache_line[k][674] = (mem_line[line_addr][674] & (~hit)) | (cache_line[k][674] & (hit));
				cache_line[k][675] = (mem_line[line_addr][675] & (~hit)) | (cache_line[k][675] & (hit));
				cache_line[k][676] = (mem_line[line_addr][676] & (~hit)) | (cache_line[k][676] & (hit));
				cache_line[k][677] = (mem_line[line_addr][677] & (~hit)) | (cache_line[k][677] & (hit));
				cache_line[k][678] = (mem_line[line_addr][678] & (~hit)) | (cache_line[k][678] & (hit));
				cache_line[k][679] = (mem_line[line_addr][679] & (~hit)) | (cache_line[k][679] & (hit));
				cache_line[k][680] = (mem_line[line_addr][680] & (~hit)) | (cache_line[k][680] & (hit));
				cache_line[k][681] = (mem_line[line_addr][681] & (~hit)) | (cache_line[k][681] & (hit));
				cache_line[k][682] = (mem_line[line_addr][682] & (~hit)) | (cache_line[k][682] & (hit));
				cache_line[k][683] = (mem_line[line_addr][683] & (~hit)) | (cache_line[k][683] & (hit));
				cache_line[k][684] = (mem_line[line_addr][684] & (~hit)) | (cache_line[k][684] & (hit));
				cache_line[k][685] = (mem_line[line_addr][685] & (~hit)) | (cache_line[k][685] & (hit));
				cache_line[k][686] = (mem_line[line_addr][686] & (~hit)) | (cache_line[k][686] & (hit));
				cache_line[k][687] = (mem_line[line_addr][687] & (~hit)) | (cache_line[k][687] & (hit));
				cache_line[k][688] = (mem_line[line_addr][688] & (~hit)) | (cache_line[k][688] & (hit));
				cache_line[k][689] = (mem_line[line_addr][689] & (~hit)) | (cache_line[k][689] & (hit));
				cache_line[k][690] = (mem_line[line_addr][690] & (~hit)) | (cache_line[k][690] & (hit));
				cache_line[k][691] = (mem_line[line_addr][691] & (~hit)) | (cache_line[k][691] & (hit));
				cache_line[k][692] = (mem_line[line_addr][692] & (~hit)) | (cache_line[k][692] & (hit));
				cache_line[k][693] = (mem_line[line_addr][693] & (~hit)) | (cache_line[k][693] & (hit));
				cache_line[k][694] = (mem_line[line_addr][694] & (~hit)) | (cache_line[k][694] & (hit));
				cache_line[k][695] = (mem_line[line_addr][695] & (~hit)) | (cache_line[k][695] & (hit));
				cache_line[k][696] = (mem_line[line_addr][696] & (~hit)) | (cache_line[k][696] & (hit));
				cache_line[k][697] = (mem_line[line_addr][697] & (~hit)) | (cache_line[k][697] & (hit));
				cache_line[k][698] = (mem_line[line_addr][698] & (~hit)) | (cache_line[k][698] & (hit));
				cache_line[k][699] = (mem_line[line_addr][699] & (~hit)) | (cache_line[k][699] & (hit));
				cache_line[k][700] = (mem_line[line_addr][700] & (~hit)) | (cache_line[k][700] & (hit));
				cache_line[k][701] = (mem_line[line_addr][701] & (~hit)) | (cache_line[k][701] & (hit));
				cache_line[k][702] = (mem_line[line_addr][702] & (~hit)) | (cache_line[k][702] & (hit));
				cache_line[k][703] = (mem_line[line_addr][703] & (~hit)) | (cache_line[k][703] & (hit));
				cache_line[k][704] = (mem_line[line_addr][704] & (~hit)) | (cache_line[k][704] & (hit));
				cache_line[k][705] = (mem_line[line_addr][705] & (~hit)) | (cache_line[k][705] & (hit));
				cache_line[k][706] = (mem_line[line_addr][706] & (~hit)) | (cache_line[k][706] & (hit));
				cache_line[k][707] = (mem_line[line_addr][707] & (~hit)) | (cache_line[k][707] & (hit));
				cache_line[k][708] = (mem_line[line_addr][708] & (~hit)) | (cache_line[k][708] & (hit));
				cache_line[k][709] = (mem_line[line_addr][709] & (~hit)) | (cache_line[k][709] & (hit));
				cache_line[k][710] = (mem_line[line_addr][710] & (~hit)) | (cache_line[k][710] & (hit));
				cache_line[k][711] = (mem_line[line_addr][711] & (~hit)) | (cache_line[k][711] & (hit));
				cache_line[k][712] = (mem_line[line_addr][712] & (~hit)) | (cache_line[k][712] & (hit));
				cache_line[k][713] = (mem_line[line_addr][713] & (~hit)) | (cache_line[k][713] & (hit));
				cache_line[k][714] = (mem_line[line_addr][714] & (~hit)) | (cache_line[k][714] & (hit));
				cache_line[k][715] = (mem_line[line_addr][715] & (~hit)) | (cache_line[k][715] & (hit));
				cache_line[k][716] = (mem_line[line_addr][716] & (~hit)) | (cache_line[k][716] & (hit));
				cache_line[k][717] = (mem_line[line_addr][717] & (~hit)) | (cache_line[k][717] & (hit));
				cache_line[k][718] = (mem_line[line_addr][718] & (~hit)) | (cache_line[k][718] & (hit));
				cache_line[k][719] = (mem_line[line_addr][719] & (~hit)) | (cache_line[k][719] & (hit));
				cache_line[k][720] = (mem_line[line_addr][720] & (~hit)) | (cache_line[k][720] & (hit));
				cache_line[k][721] = (mem_line[line_addr][721] & (~hit)) | (cache_line[k][721] & (hit));
				cache_line[k][722] = (mem_line[line_addr][722] & (~hit)) | (cache_line[k][722] & (hit));
				cache_line[k][723] = (mem_line[line_addr][723] & (~hit)) | (cache_line[k][723] & (hit));
				cache_line[k][724] = (mem_line[line_addr][724] & (~hit)) | (cache_line[k][724] & (hit));
				cache_line[k][725] = (mem_line[line_addr][725] & (~hit)) | (cache_line[k][725] & (hit));
				cache_line[k][726] = (mem_line[line_addr][726] & (~hit)) | (cache_line[k][726] & (hit));
				cache_line[k][727] = (mem_line[line_addr][727] & (~hit)) | (cache_line[k][727] & (hit));
				cache_line[k][728] = (mem_line[line_addr][728] & (~hit)) | (cache_line[k][728] & (hit));
				cache_line[k][729] = (mem_line[line_addr][729] & (~hit)) | (cache_line[k][729] & (hit));
				cache_line[k][730] = (mem_line[line_addr][730] & (~hit)) | (cache_line[k][730] & (hit));
				cache_line[k][731] = (mem_line[line_addr][731] & (~hit)) | (cache_line[k][731] & (hit));
				cache_line[k][732] = (mem_line[line_addr][732] & (~hit)) | (cache_line[k][732] & (hit));
				cache_line[k][733] = (mem_line[line_addr][733] & (~hit)) | (cache_line[k][733] & (hit));
				cache_line[k][734] = (mem_line[line_addr][734] & (~hit)) | (cache_line[k][734] & (hit));
				cache_line[k][735] = (mem_line[line_addr][735] & (~hit)) | (cache_line[k][735] & (hit));
				cache_line[k][736] = (mem_line[line_addr][736] & (~hit)) | (cache_line[k][736] & (hit));
				cache_line[k][737] = (mem_line[line_addr][737] & (~hit)) | (cache_line[k][737] & (hit));
				cache_line[k][738] = (mem_line[line_addr][738] & (~hit)) | (cache_line[k][738] & (hit));
				cache_line[k][739] = (mem_line[line_addr][739] & (~hit)) | (cache_line[k][739] & (hit));
				cache_line[k][740] = (mem_line[line_addr][740] & (~hit)) | (cache_line[k][740] & (hit));
				cache_line[k][741] = (mem_line[line_addr][741] & (~hit)) | (cache_line[k][741] & (hit));
				cache_line[k][742] = (mem_line[line_addr][742] & (~hit)) | (cache_line[k][742] & (hit));
				cache_line[k][743] = (mem_line[line_addr][743] & (~hit)) | (cache_line[k][743] & (hit));
				cache_line[k][744] = (mem_line[line_addr][744] & (~hit)) | (cache_line[k][744] & (hit));
				cache_line[k][745] = (mem_line[line_addr][745] & (~hit)) | (cache_line[k][745] & (hit));
				cache_line[k][746] = (mem_line[line_addr][746] & (~hit)) | (cache_line[k][746] & (hit));
				cache_line[k][747] = (mem_line[line_addr][747] & (~hit)) | (cache_line[k][747] & (hit));
				cache_line[k][748] = (mem_line[line_addr][748] & (~hit)) | (cache_line[k][748] & (hit));
				cache_line[k][749] = (mem_line[line_addr][749] & (~hit)) | (cache_line[k][749] & (hit));
				cache_line[k][750] = (mem_line[line_addr][750] & (~hit)) | (cache_line[k][750] & (hit));
				cache_line[k][751] = (mem_line[line_addr][751] & (~hit)) | (cache_line[k][751] & (hit));
				cache_line[k][752] = (mem_line[line_addr][752] & (~hit)) | (cache_line[k][752] & (hit));
				cache_line[k][753] = (mem_line[line_addr][753] & (~hit)) | (cache_line[k][753] & (hit));
				cache_line[k][754] = (mem_line[line_addr][754] & (~hit)) | (cache_line[k][754] & (hit));
				cache_line[k][755] = (mem_line[line_addr][755] & (~hit)) | (cache_line[k][755] & (hit));
				cache_line[k][756] = (mem_line[line_addr][756] & (~hit)) | (cache_line[k][756] & (hit));
				cache_line[k][757] = (mem_line[line_addr][757] & (~hit)) | (cache_line[k][757] & (hit));
				cache_line[k][758] = (mem_line[line_addr][758] & (~hit)) | (cache_line[k][758] & (hit));
				cache_line[k][759] = (mem_line[line_addr][759] & (~hit)) | (cache_line[k][759] & (hit));
				cache_line[k][760] = (mem_line[line_addr][760] & (~hit)) | (cache_line[k][760] & (hit));
				cache_line[k][761] = (mem_line[line_addr][761] & (~hit)) | (cache_line[k][761] & (hit));
				cache_line[k][762] = (mem_line[line_addr][762] & (~hit)) | (cache_line[k][762] & (hit));
				cache_line[k][763] = (mem_line[line_addr][763] & (~hit)) | (cache_line[k][763] & (hit));
				cache_line[k][764] = (mem_line[line_addr][764] & (~hit)) | (cache_line[k][764] & (hit));
				cache_line[k][765] = (mem_line[line_addr][765] & (~hit)) | (cache_line[k][765] & (hit));
				cache_line[k][766] = (mem_line[line_addr][766] & (~hit)) | (cache_line[k][766] & (hit));
				cache_line[k][767] = (mem_line[line_addr][767] & (~hit)) | (cache_line[k][767] & (hit));
				cache_line[k][768] = (mem_line[line_addr][768] & (~hit)) | (cache_line[k][768] & (hit));
				cache_line[k][769] = (mem_line[line_addr][769] & (~hit)) | (cache_line[k][769] & (hit));
				cache_line[k][770] = (mem_line[line_addr][770] & (~hit)) | (cache_line[k][770] & (hit));
				cache_line[k][771] = (mem_line[line_addr][771] & (~hit)) | (cache_line[k][771] & (hit));
				cache_line[k][772] = (mem_line[line_addr][772] & (~hit)) | (cache_line[k][772] & (hit));
				cache_line[k][773] = (mem_line[line_addr][773] & (~hit)) | (cache_line[k][773] & (hit));
				cache_line[k][774] = (mem_line[line_addr][774] & (~hit)) | (cache_line[k][774] & (hit));
				cache_line[k][775] = (mem_line[line_addr][775] & (~hit)) | (cache_line[k][775] & (hit));
				cache_line[k][776] = (mem_line[line_addr][776] & (~hit)) | (cache_line[k][776] & (hit));
				cache_line[k][777] = (mem_line[line_addr][777] & (~hit)) | (cache_line[k][777] & (hit));
				cache_line[k][778] = (mem_line[line_addr][778] & (~hit)) | (cache_line[k][778] & (hit));
				cache_line[k][779] = (mem_line[line_addr][779] & (~hit)) | (cache_line[k][779] & (hit));
				cache_line[k][780] = (mem_line[line_addr][780] & (~hit)) | (cache_line[k][780] & (hit));
				cache_line[k][781] = (mem_line[line_addr][781] & (~hit)) | (cache_line[k][781] & (hit));
				cache_line[k][782] = (mem_line[line_addr][782] & (~hit)) | (cache_line[k][782] & (hit));
				cache_line[k][783] = (mem_line[line_addr][783] & (~hit)) | (cache_line[k][783] & (hit));
				cache_line[k][784] = (mem_line[line_addr][784] & (~hit)) | (cache_line[k][784] & (hit));
				cache_line[k][785] = (mem_line[line_addr][785] & (~hit)) | (cache_line[k][785] & (hit));
				cache_line[k][786] = (mem_line[line_addr][786] & (~hit)) | (cache_line[k][786] & (hit));
				cache_line[k][787] = (mem_line[line_addr][787] & (~hit)) | (cache_line[k][787] & (hit));
				cache_line[k][788] = (mem_line[line_addr][788] & (~hit)) | (cache_line[k][788] & (hit));
				cache_line[k][789] = (mem_line[line_addr][789] & (~hit)) | (cache_line[k][789] & (hit));
				cache_line[k][790] = (mem_line[line_addr][790] & (~hit)) | (cache_line[k][790] & (hit));
				cache_line[k][791] = (mem_line[line_addr][791] & (~hit)) | (cache_line[k][791] & (hit));
				cache_line[k][792] = (mem_line[line_addr][792] & (~hit)) | (cache_line[k][792] & (hit));
				cache_line[k][793] = (mem_line[line_addr][793] & (~hit)) | (cache_line[k][793] & (hit));
				cache_line[k][794] = (mem_line[line_addr][794] & (~hit)) | (cache_line[k][794] & (hit));
				cache_line[k][795] = (mem_line[line_addr][795] & (~hit)) | (cache_line[k][795] & (hit));
				cache_line[k][796] = (mem_line[line_addr][796] & (~hit)) | (cache_line[k][796] & (hit));
				cache_line[k][797] = (mem_line[line_addr][797] & (~hit)) | (cache_line[k][797] & (hit));
				cache_line[k][798] = (mem_line[line_addr][798] & (~hit)) | (cache_line[k][798] & (hit));
				cache_line[k][799] = (mem_line[line_addr][799] & (~hit)) | (cache_line[k][799] & (hit));
				cache_line[k][800] = (mem_line[line_addr][800] & (~hit)) | (cache_line[k][800] & (hit));
				cache_line[k][801] = (mem_line[line_addr][801] & (~hit)) | (cache_line[k][801] & (hit));
				cache_line[k][802] = (mem_line[line_addr][802] & (~hit)) | (cache_line[k][802] & (hit));
				cache_line[k][803] = (mem_line[line_addr][803] & (~hit)) | (cache_line[k][803] & (hit));
				cache_line[k][804] = (mem_line[line_addr][804] & (~hit)) | (cache_line[k][804] & (hit));
				cache_line[k][805] = (mem_line[line_addr][805] & (~hit)) | (cache_line[k][805] & (hit));
				cache_line[k][806] = (mem_line[line_addr][806] & (~hit)) | (cache_line[k][806] & (hit));
				cache_line[k][807] = (mem_line[line_addr][807] & (~hit)) | (cache_line[k][807] & (hit));
				cache_line[k][808] = (mem_line[line_addr][808] & (~hit)) | (cache_line[k][808] & (hit));
				cache_line[k][809] = (mem_line[line_addr][809] & (~hit)) | (cache_line[k][809] & (hit));
				cache_line[k][810] = (mem_line[line_addr][810] & (~hit)) | (cache_line[k][810] & (hit));
				cache_line[k][811] = (mem_line[line_addr][811] & (~hit)) | (cache_line[k][811] & (hit));
				cache_line[k][812] = (mem_line[line_addr][812] & (~hit)) | (cache_line[k][812] & (hit));
				cache_line[k][813] = (mem_line[line_addr][813] & (~hit)) | (cache_line[k][813] & (hit));
				cache_line[k][814] = (mem_line[line_addr][814] & (~hit)) | (cache_line[k][814] & (hit));
				cache_line[k][815] = (mem_line[line_addr][815] & (~hit)) | (cache_line[k][815] & (hit));
				cache_line[k][816] = (mem_line[line_addr][816] & (~hit)) | (cache_line[k][816] & (hit));
				cache_line[k][817] = (mem_line[line_addr][817] & (~hit)) | (cache_line[k][817] & (hit));
				cache_line[k][818] = (mem_line[line_addr][818] & (~hit)) | (cache_line[k][818] & (hit));
				cache_line[k][819] = (mem_line[line_addr][819] & (~hit)) | (cache_line[k][819] & (hit));
				cache_line[k][820] = (mem_line[line_addr][820] & (~hit)) | (cache_line[k][820] & (hit));
				cache_line[k][821] = (mem_line[line_addr][821] & (~hit)) | (cache_line[k][821] & (hit));
				cache_line[k][822] = (mem_line[line_addr][822] & (~hit)) | (cache_line[k][822] & (hit));
				cache_line[k][823] = (mem_line[line_addr][823] & (~hit)) | (cache_line[k][823] & (hit));
				cache_line[k][824] = (mem_line[line_addr][824] & (~hit)) | (cache_line[k][824] & (hit));
				cache_line[k][825] = (mem_line[line_addr][825] & (~hit)) | (cache_line[k][825] & (hit));
				cache_line[k][826] = (mem_line[line_addr][826] & (~hit)) | (cache_line[k][826] & (hit));
				cache_line[k][827] = (mem_line[line_addr][827] & (~hit)) | (cache_line[k][827] & (hit));
				cache_line[k][828] = (mem_line[line_addr][828] & (~hit)) | (cache_line[k][828] & (hit));
				cache_line[k][829] = (mem_line[line_addr][829] & (~hit)) | (cache_line[k][829] & (hit));
				cache_line[k][830] = (mem_line[line_addr][830] & (~hit)) | (cache_line[k][830] & (hit));
				cache_line[k][831] = (mem_line[line_addr][831] & (~hit)) | (cache_line[k][831] & (hit));
				cache_line[k][832] = (mem_line[line_addr][832] & (~hit)) | (cache_line[k][832] & (hit));
				cache_line[k][833] = (mem_line[line_addr][833] & (~hit)) | (cache_line[k][833] & (hit));
				cache_line[k][834] = (mem_line[line_addr][834] & (~hit)) | (cache_line[k][834] & (hit));
				cache_line[k][835] = (mem_line[line_addr][835] & (~hit)) | (cache_line[k][835] & (hit));
				cache_line[k][836] = (mem_line[line_addr][836] & (~hit)) | (cache_line[k][836] & (hit));
				cache_line[k][837] = (mem_line[line_addr][837] & (~hit)) | (cache_line[k][837] & (hit));
				cache_line[k][838] = (mem_line[line_addr][838] & (~hit)) | (cache_line[k][838] & (hit));
				cache_line[k][839] = (mem_line[line_addr][839] & (~hit)) | (cache_line[k][839] & (hit));
				cache_line[k][840] = (mem_line[line_addr][840] & (~hit)) | (cache_line[k][840] & (hit));
				cache_line[k][841] = (mem_line[line_addr][841] & (~hit)) | (cache_line[k][841] & (hit));
				cache_line[k][842] = (mem_line[line_addr][842] & (~hit)) | (cache_line[k][842] & (hit));
				cache_line[k][843] = (mem_line[line_addr][843] & (~hit)) | (cache_line[k][843] & (hit));
				cache_line[k][844] = (mem_line[line_addr][844] & (~hit)) | (cache_line[k][844] & (hit));
				cache_line[k][845] = (mem_line[line_addr][845] & (~hit)) | (cache_line[k][845] & (hit));
				cache_line[k][846] = (mem_line[line_addr][846] & (~hit)) | (cache_line[k][846] & (hit));
				cache_line[k][847] = (mem_line[line_addr][847] & (~hit)) | (cache_line[k][847] & (hit));
				cache_line[k][848] = (mem_line[line_addr][848] & (~hit)) | (cache_line[k][848] & (hit));
				cache_line[k][849] = (mem_line[line_addr][849] & (~hit)) | (cache_line[k][849] & (hit));
				cache_line[k][850] = (mem_line[line_addr][850] & (~hit)) | (cache_line[k][850] & (hit));
				cache_line[k][851] = (mem_line[line_addr][851] & (~hit)) | (cache_line[k][851] & (hit));
				cache_line[k][852] = (mem_line[line_addr][852] & (~hit)) | (cache_line[k][852] & (hit));
				cache_line[k][853] = (mem_line[line_addr][853] & (~hit)) | (cache_line[k][853] & (hit));
				cache_line[k][854] = (mem_line[line_addr][854] & (~hit)) | (cache_line[k][854] & (hit));
				cache_line[k][855] = (mem_line[line_addr][855] & (~hit)) | (cache_line[k][855] & (hit));
				cache_line[k][856] = (mem_line[line_addr][856] & (~hit)) | (cache_line[k][856] & (hit));
				cache_line[k][857] = (mem_line[line_addr][857] & (~hit)) | (cache_line[k][857] & (hit));
				cache_line[k][858] = (mem_line[line_addr][858] & (~hit)) | (cache_line[k][858] & (hit));
				cache_line[k][859] = (mem_line[line_addr][859] & (~hit)) | (cache_line[k][859] & (hit));
				cache_line[k][860] = (mem_line[line_addr][860] & (~hit)) | (cache_line[k][860] & (hit));
				cache_line[k][861] = (mem_line[line_addr][861] & (~hit)) | (cache_line[k][861] & (hit));
				cache_line[k][862] = (mem_line[line_addr][862] & (~hit)) | (cache_line[k][862] & (hit));
				cache_line[k][863] = (mem_line[line_addr][863] & (~hit)) | (cache_line[k][863] & (hit));
				cache_line[k][864] = (mem_line[line_addr][864] & (~hit)) | (cache_line[k][864] & (hit));
				cache_line[k][865] = (mem_line[line_addr][865] & (~hit)) | (cache_line[k][865] & (hit));
				cache_line[k][866] = (mem_line[line_addr][866] & (~hit)) | (cache_line[k][866] & (hit));
				cache_line[k][867] = (mem_line[line_addr][867] & (~hit)) | (cache_line[k][867] & (hit));
				cache_line[k][868] = (mem_line[line_addr][868] & (~hit)) | (cache_line[k][868] & (hit));
				cache_line[k][869] = (mem_line[line_addr][869] & (~hit)) | (cache_line[k][869] & (hit));
				cache_line[k][870] = (mem_line[line_addr][870] & (~hit)) | (cache_line[k][870] & (hit));
				cache_line[k][871] = (mem_line[line_addr][871] & (~hit)) | (cache_line[k][871] & (hit));
				cache_line[k][872] = (mem_line[line_addr][872] & (~hit)) | (cache_line[k][872] & (hit));
				cache_line[k][873] = (mem_line[line_addr][873] & (~hit)) | (cache_line[k][873] & (hit));
				cache_line[k][874] = (mem_line[line_addr][874] & (~hit)) | (cache_line[k][874] & (hit));
				cache_line[k][875] = (mem_line[line_addr][875] & (~hit)) | (cache_line[k][875] & (hit));
				cache_line[k][876] = (mem_line[line_addr][876] & (~hit)) | (cache_line[k][876] & (hit));
				cache_line[k][877] = (mem_line[line_addr][877] & (~hit)) | (cache_line[k][877] & (hit));
				cache_line[k][878] = (mem_line[line_addr][878] & (~hit)) | (cache_line[k][878] & (hit));
				cache_line[k][879] = (mem_line[line_addr][879] & (~hit)) | (cache_line[k][879] & (hit));
				cache_line[k][880] = (mem_line[line_addr][880] & (~hit)) | (cache_line[k][880] & (hit));
				cache_line[k][881] = (mem_line[line_addr][881] & (~hit)) | (cache_line[k][881] & (hit));
				cache_line[k][882] = (mem_line[line_addr][882] & (~hit)) | (cache_line[k][882] & (hit));
				cache_line[k][883] = (mem_line[line_addr][883] & (~hit)) | (cache_line[k][883] & (hit));
				cache_line[k][884] = (mem_line[line_addr][884] & (~hit)) | (cache_line[k][884] & (hit));
				cache_line[k][885] = (mem_line[line_addr][885] & (~hit)) | (cache_line[k][885] & (hit));
				cache_line[k][886] = (mem_line[line_addr][886] & (~hit)) | (cache_line[k][886] & (hit));
				cache_line[k][887] = (mem_line[line_addr][887] & (~hit)) | (cache_line[k][887] & (hit));
				cache_line[k][888] = (mem_line[line_addr][888] & (~hit)) | (cache_line[k][888] & (hit));
				cache_line[k][889] = (mem_line[line_addr][889] & (~hit)) | (cache_line[k][889] & (hit));
				cache_line[k][890] = (mem_line[line_addr][890] & (~hit)) | (cache_line[k][890] & (hit));
				cache_line[k][891] = (mem_line[line_addr][891] & (~hit)) | (cache_line[k][891] & (hit));
				cache_line[k][892] = (mem_line[line_addr][892] & (~hit)) | (cache_line[k][892] & (hit));
				cache_line[k][893] = (mem_line[line_addr][893] & (~hit)) | (cache_line[k][893] & (hit));
				cache_line[k][894] = (mem_line[line_addr][894] & (~hit)) | (cache_line[k][894] & (hit));
				cache_line[k][895] = (mem_line[line_addr][895] & (~hit)) | (cache_line[k][895] & (hit));
				cache_line[k][896] = (mem_line[line_addr][896] & (~hit)) | (cache_line[k][896] & (hit));
				cache_line[k][897] = (mem_line[line_addr][897] & (~hit)) | (cache_line[k][897] & (hit));
				cache_line[k][898] = (mem_line[line_addr][898] & (~hit)) | (cache_line[k][898] & (hit));
				cache_line[k][899] = (mem_line[line_addr][899] & (~hit)) | (cache_line[k][899] & (hit));
				cache_line[k][900] = (mem_line[line_addr][900] & (~hit)) | (cache_line[k][900] & (hit));
				cache_line[k][901] = (mem_line[line_addr][901] & (~hit)) | (cache_line[k][901] & (hit));
				cache_line[k][902] = (mem_line[line_addr][902] & (~hit)) | (cache_line[k][902] & (hit));
				cache_line[k][903] = (mem_line[line_addr][903] & (~hit)) | (cache_line[k][903] & (hit));
				cache_line[k][904] = (mem_line[line_addr][904] & (~hit)) | (cache_line[k][904] & (hit));
				cache_line[k][905] = (mem_line[line_addr][905] & (~hit)) | (cache_line[k][905] & (hit));
				cache_line[k][906] = (mem_line[line_addr][906] & (~hit)) | (cache_line[k][906] & (hit));
				cache_line[k][907] = (mem_line[line_addr][907] & (~hit)) | (cache_line[k][907] & (hit));
				cache_line[k][908] = (mem_line[line_addr][908] & (~hit)) | (cache_line[k][908] & (hit));
				cache_line[k][909] = (mem_line[line_addr][909] & (~hit)) | (cache_line[k][909] & (hit));
				cache_line[k][910] = (mem_line[line_addr][910] & (~hit)) | (cache_line[k][910] & (hit));
				cache_line[k][911] = (mem_line[line_addr][911] & (~hit)) | (cache_line[k][911] & (hit));
				cache_line[k][912] = (mem_line[line_addr][912] & (~hit)) | (cache_line[k][912] & (hit));
				cache_line[k][913] = (mem_line[line_addr][913] & (~hit)) | (cache_line[k][913] & (hit));
				cache_line[k][914] = (mem_line[line_addr][914] & (~hit)) | (cache_line[k][914] & (hit));
				cache_line[k][915] = (mem_line[line_addr][915] & (~hit)) | (cache_line[k][915] & (hit));
				cache_line[k][916] = (mem_line[line_addr][916] & (~hit)) | (cache_line[k][916] & (hit));
				cache_line[k][917] = (mem_line[line_addr][917] & (~hit)) | (cache_line[k][917] & (hit));
				cache_line[k][918] = (mem_line[line_addr][918] & (~hit)) | (cache_line[k][918] & (hit));
				cache_line[k][919] = (mem_line[line_addr][919] & (~hit)) | (cache_line[k][919] & (hit));
				cache_line[k][920] = (mem_line[line_addr][920] & (~hit)) | (cache_line[k][920] & (hit));
				cache_line[k][921] = (mem_line[line_addr][921] & (~hit)) | (cache_line[k][921] & (hit));
				cache_line[k][922] = (mem_line[line_addr][922] & (~hit)) | (cache_line[k][922] & (hit));
				cache_line[k][923] = (mem_line[line_addr][923] & (~hit)) | (cache_line[k][923] & (hit));
				cache_line[k][924] = (mem_line[line_addr][924] & (~hit)) | (cache_line[k][924] & (hit));
				cache_line[k][925] = (mem_line[line_addr][925] & (~hit)) | (cache_line[k][925] & (hit));
				cache_line[k][926] = (mem_line[line_addr][926] & (~hit)) | (cache_line[k][926] & (hit));
				cache_line[k][927] = (mem_line[line_addr][927] & (~hit)) | (cache_line[k][927] & (hit));
				cache_line[k][928] = (mem_line[line_addr][928] & (~hit)) | (cache_line[k][928] & (hit));
				cache_line[k][929] = (mem_line[line_addr][929] & (~hit)) | (cache_line[k][929] & (hit));
				cache_line[k][930] = (mem_line[line_addr][930] & (~hit)) | (cache_line[k][930] & (hit));
				cache_line[k][931] = (mem_line[line_addr][931] & (~hit)) | (cache_line[k][931] & (hit));
				cache_line[k][932] = (mem_line[line_addr][932] & (~hit)) | (cache_line[k][932] & (hit));
				cache_line[k][933] = (mem_line[line_addr][933] & (~hit)) | (cache_line[k][933] & (hit));
				cache_line[k][934] = (mem_line[line_addr][934] & (~hit)) | (cache_line[k][934] & (hit));
				cache_line[k][935] = (mem_line[line_addr][935] & (~hit)) | (cache_line[k][935] & (hit));
				cache_line[k][936] = (mem_line[line_addr][936] & (~hit)) | (cache_line[k][936] & (hit));
				cache_line[k][937] = (mem_line[line_addr][937] & (~hit)) | (cache_line[k][937] & (hit));
				cache_line[k][938] = (mem_line[line_addr][938] & (~hit)) | (cache_line[k][938] & (hit));
				cache_line[k][939] = (mem_line[line_addr][939] & (~hit)) | (cache_line[k][939] & (hit));
				cache_line[k][940] = (mem_line[line_addr][940] & (~hit)) | (cache_line[k][940] & (hit));
				cache_line[k][941] = (mem_line[line_addr][941] & (~hit)) | (cache_line[k][941] & (hit));
				cache_line[k][942] = (mem_line[line_addr][942] & (~hit)) | (cache_line[k][942] & (hit));
				cache_line[k][943] = (mem_line[line_addr][943] & (~hit)) | (cache_line[k][943] & (hit));
				cache_line[k][944] = (mem_line[line_addr][944] & (~hit)) | (cache_line[k][944] & (hit));
				cache_line[k][945] = (mem_line[line_addr][945] & (~hit)) | (cache_line[k][945] & (hit));
				cache_line[k][946] = (mem_line[line_addr][946] & (~hit)) | (cache_line[k][946] & (hit));
				cache_line[k][947] = (mem_line[line_addr][947] & (~hit)) | (cache_line[k][947] & (hit));
				cache_line[k][948] = (mem_line[line_addr][948] & (~hit)) | (cache_line[k][948] & (hit));
				cache_line[k][949] = (mem_line[line_addr][949] & (~hit)) | (cache_line[k][949] & (hit));
				cache_line[k][950] = (mem_line[line_addr][950] & (~hit)) | (cache_line[k][950] & (hit));
				cache_line[k][951] = (mem_line[line_addr][951] & (~hit)) | (cache_line[k][951] & (hit));
				cache_line[k][952] = (mem_line[line_addr][952] & (~hit)) | (cache_line[k][952] & (hit));
				cache_line[k][953] = (mem_line[line_addr][953] & (~hit)) | (cache_line[k][953] & (hit));
				cache_line[k][954] = (mem_line[line_addr][954] & (~hit)) | (cache_line[k][954] & (hit));
				cache_line[k][955] = (mem_line[line_addr][955] & (~hit)) | (cache_line[k][955] & (hit));
				cache_line[k][956] = (mem_line[line_addr][956] & (~hit)) | (cache_line[k][956] & (hit));
				cache_line[k][957] = (mem_line[line_addr][957] & (~hit)) | (cache_line[k][957] & (hit));
				cache_line[k][958] = (mem_line[line_addr][958] & (~hit)) | (cache_line[k][958] & (hit));
				cache_line[k][959] = (mem_line[line_addr][959] & (~hit)) | (cache_line[k][959] & (hit));
				cache_line[k][960] = (mem_line[line_addr][960] & (~hit)) | (cache_line[k][960] & (hit));
				cache_line[k][961] = (mem_line[line_addr][961] & (~hit)) | (cache_line[k][961] & (hit));
				cache_line[k][962] = (mem_line[line_addr][962] & (~hit)) | (cache_line[k][962] & (hit));
				cache_line[k][963] = (mem_line[line_addr][963] & (~hit)) | (cache_line[k][963] & (hit));
				cache_line[k][964] = (mem_line[line_addr][964] & (~hit)) | (cache_line[k][964] & (hit));
				cache_line[k][965] = (mem_line[line_addr][965] & (~hit)) | (cache_line[k][965] & (hit));
				cache_line[k][966] = (mem_line[line_addr][966] & (~hit)) | (cache_line[k][966] & (hit));
				cache_line[k][967] = (mem_line[line_addr][967] & (~hit)) | (cache_line[k][967] & (hit));
				cache_line[k][968] = (mem_line[line_addr][968] & (~hit)) | (cache_line[k][968] & (hit));
				cache_line[k][969] = (mem_line[line_addr][969] & (~hit)) | (cache_line[k][969] & (hit));
				cache_line[k][970] = (mem_line[line_addr][970] & (~hit)) | (cache_line[k][970] & (hit));
				cache_line[k][971] = (mem_line[line_addr][971] & (~hit)) | (cache_line[k][971] & (hit));
				cache_line[k][972] = (mem_line[line_addr][972] & (~hit)) | (cache_line[k][972] & (hit));
				cache_line[k][973] = (mem_line[line_addr][973] & (~hit)) | (cache_line[k][973] & (hit));
				cache_line[k][974] = (mem_line[line_addr][974] & (~hit)) | (cache_line[k][974] & (hit));
				cache_line[k][975] = (mem_line[line_addr][975] & (~hit)) | (cache_line[k][975] & (hit));
				cache_line[k][976] = (mem_line[line_addr][976] & (~hit)) | (cache_line[k][976] & (hit));
				cache_line[k][977] = (mem_line[line_addr][977] & (~hit)) | (cache_line[k][977] & (hit));
				cache_line[k][978] = (mem_line[line_addr][978] & (~hit)) | (cache_line[k][978] & (hit));
				cache_line[k][979] = (mem_line[line_addr][979] & (~hit)) | (cache_line[k][979] & (hit));
				cache_line[k][980] = (mem_line[line_addr][980] & (~hit)) | (cache_line[k][980] & (hit));
				cache_line[k][981] = (mem_line[line_addr][981] & (~hit)) | (cache_line[k][981] & (hit));
				cache_line[k][982] = (mem_line[line_addr][982] & (~hit)) | (cache_line[k][982] & (hit));
				cache_line[k][983] = (mem_line[line_addr][983] & (~hit)) | (cache_line[k][983] & (hit));
				cache_line[k][984] = (mem_line[line_addr][984] & (~hit)) | (cache_line[k][984] & (hit));
				cache_line[k][985] = (mem_line[line_addr][985] & (~hit)) | (cache_line[k][985] & (hit));
				cache_line[k][986] = (mem_line[line_addr][986] & (~hit)) | (cache_line[k][986] & (hit));
				cache_line[k][987] = (mem_line[line_addr][987] & (~hit)) | (cache_line[k][987] & (hit));
				cache_line[k][988] = (mem_line[line_addr][988] & (~hit)) | (cache_line[k][988] & (hit));
				cache_line[k][989] = (mem_line[line_addr][989] & (~hit)) | (cache_line[k][989] & (hit));
				cache_line[k][990] = (mem_line[line_addr][990] & (~hit)) | (cache_line[k][990] & (hit));
				cache_line[k][991] = (mem_line[line_addr][991] & (~hit)) | (cache_line[k][991] & (hit));
				cache_line[k][992] = (mem_line[line_addr][992] & (~hit)) | (cache_line[k][992] & (hit));
				cache_line[k][993] = (mem_line[line_addr][993] & (~hit)) | (cache_line[k][993] & (hit));
				cache_line[k][994] = (mem_line[line_addr][994] & (~hit)) | (cache_line[k][994] & (hit));
				cache_line[k][995] = (mem_line[line_addr][995] & (~hit)) | (cache_line[k][995] & (hit));
				cache_line[k][996] = (mem_line[line_addr][996] & (~hit)) | (cache_line[k][996] & (hit));
				cache_line[k][997] = (mem_line[line_addr][997] & (~hit)) | (cache_line[k][997] & (hit));
				cache_line[k][998] = (mem_line[line_addr][998] & (~hit)) | (cache_line[k][998] & (hit));
				cache_line[k][999] = (mem_line[line_addr][999] & (~hit)) | (cache_line[k][999] & (hit));
				cache_line[k][1000] = (mem_line[line_addr][1000] & (~hit)) | (cache_line[k][1000] & (hit));
				cache_line[k][1001] = (mem_line[line_addr][1001] & (~hit)) | (cache_line[k][1001] & (hit));
				cache_line[k][1002] = (mem_line[line_addr][1002] & (~hit)) | (cache_line[k][1002] & (hit));
				cache_line[k][1003] = (mem_line[line_addr][1003] & (~hit)) | (cache_line[k][1003] & (hit));
				cache_line[k][1004] = (mem_line[line_addr][1004] & (~hit)) | (cache_line[k][1004] & (hit));
				cache_line[k][1005] = (mem_line[line_addr][1005] & (~hit)) | (cache_line[k][1005] & (hit));
				cache_line[k][1006] = (mem_line[line_addr][1006] & (~hit)) | (cache_line[k][1006] & (hit));
				cache_line[k][1007] = (mem_line[line_addr][1007] & (~hit)) | (cache_line[k][1007] & (hit));
				cache_line[k][1008] = (mem_line[line_addr][1008] & (~hit)) | (cache_line[k][1008] & (hit));
				cache_line[k][1009] = (mem_line[line_addr][1009] & (~hit)) | (cache_line[k][1009] & (hit));
				cache_line[k][1010] = (mem_line[line_addr][1010] & (~hit)) | (cache_line[k][1010] & (hit));
				cache_line[k][1011] = (mem_line[line_addr][1011] & (~hit)) | (cache_line[k][1011] & (hit));
				cache_line[k][1012] = (mem_line[line_addr][1012] & (~hit)) | (cache_line[k][1012] & (hit));
				cache_line[k][1013] = (mem_line[line_addr][1013] & (~hit)) | (cache_line[k][1013] & (hit));
				cache_line[k][1014] = (mem_line[line_addr][1014] & (~hit)) | (cache_line[k][1014] & (hit));
				cache_line[k][1015] = (mem_line[line_addr][1015] & (~hit)) | (cache_line[k][1015] & (hit));
				cache_line[k][1016] = (mem_line[line_addr][1016] & (~hit)) | (cache_line[k][1016] & (hit));
				cache_line[k][1017] = (mem_line[line_addr][1017] & (~hit)) | (cache_line[k][1017] & (hit));
				cache_line[k][1018] = (mem_line[line_addr][1018] & (~hit)) | (cache_line[k][1018] & (hit));
				cache_line[k][1019] = (mem_line[line_addr][1019] & (~hit)) | (cache_line[k][1019] & (hit));
				cache_line[k][1020] = (mem_line[line_addr][1020] & (~hit)) | (cache_line[k][1020] & (hit));
				cache_line[k][1021] = (mem_line[line_addr][1021] & (~hit)) | (cache_line[k][1021] & (hit));
				cache_line[k][1022] = (mem_line[line_addr][1022] & (~hit)) | (cache_line[k][1022] & (hit));
				cache_line[k][1023] = (mem_line[line_addr][1023] & (~hit)) | (cache_line[k][1023] & (hit));
				cache_line[k][1024] = (mem_line[line_addr][1024] & (~hit)) | (cache_line[k][1024] & (hit));
				cache_line[k][1025] = (mem_line[line_addr][1025] & (~hit)) | (cache_line[k][1025] & (hit));
				cache_line[k][1026] = (mem_line[line_addr][1026] & (~hit)) | (cache_line[k][1026] & (hit));
				cache_line[k][1027] = (mem_line[line_addr][1027] & (~hit)) | (cache_line[k][1027] & (hit));
				cache_line[k][1028] = (mem_line[line_addr][1028] & (~hit)) | (cache_line[k][1028] & (hit));
				cache_line[k][1029] = (mem_line[line_addr][1029] & (~hit)) | (cache_line[k][1029] & (hit));
				cache_line[k][1030] = (mem_line[line_addr][1030] & (~hit)) | (cache_line[k][1030] & (hit));
				cache_line[k][1031] = (mem_line[line_addr][1031] & (~hit)) | (cache_line[k][1031] & (hit));
				cache_line[k][1032] = (mem_line[line_addr][1032] & (~hit)) | (cache_line[k][1032] & (hit));
				cache_line[k][1033] = (mem_line[line_addr][1033] & (~hit)) | (cache_line[k][1033] & (hit));
				cache_line[k][1034] = (mem_line[line_addr][1034] & (~hit)) | (cache_line[k][1034] & (hit));
				cache_line[k][1035] = (mem_line[line_addr][1035] & (~hit)) | (cache_line[k][1035] & (hit));
				cache_line[k][1036] = (mem_line[line_addr][1036] & (~hit)) | (cache_line[k][1036] & (hit));
				cache_line[k][1037] = (mem_line[line_addr][1037] & (~hit)) | (cache_line[k][1037] & (hit));
				cache_line[k][1038] = (mem_line[line_addr][1038] & (~hit)) | (cache_line[k][1038] & (hit));
				cache_line[k][1039] = (mem_line[line_addr][1039] & (~hit)) | (cache_line[k][1039] & (hit));
				cache_line[k][1040] = (mem_line[line_addr][1040] & (~hit)) | (cache_line[k][1040] & (hit));
				cache_line[k][1041] = (mem_line[line_addr][1041] & (~hit)) | (cache_line[k][1041] & (hit));
				cache_line[k][1042] = (mem_line[line_addr][1042] & (~hit)) | (cache_line[k][1042] & (hit));
				cache_line[k][1043] = (mem_line[line_addr][1043] & (~hit)) | (cache_line[k][1043] & (hit));
				cache_line[k][1044] = (mem_line[line_addr][1044] & (~hit)) | (cache_line[k][1044] & (hit));
				cache_line[k][1045] = (mem_line[line_addr][1045] & (~hit)) | (cache_line[k][1045] & (hit));
				cache_line[k][1046] = (mem_line[line_addr][1046] & (~hit)) | (cache_line[k][1046] & (hit));
				cache_line[k][1047] = (mem_line[line_addr][1047] & (~hit)) | (cache_line[k][1047] & (hit));
				cache_line[k][1048] = (mem_line[line_addr][1048] & (~hit)) | (cache_line[k][1048] & (hit));
				cache_line[k][1049] = (mem_line[line_addr][1049] & (~hit)) | (cache_line[k][1049] & (hit));
				cache_line[k][1050] = (mem_line[line_addr][1050] & (~hit)) | (cache_line[k][1050] & (hit));
				cache_line[k][1051] = (mem_line[line_addr][1051] & (~hit)) | (cache_line[k][1051] & (hit));
				cache_line[k][1052] = (mem_line[line_addr][1052] & (~hit)) | (cache_line[k][1052] & (hit));
				cache_line[k][1053] = (mem_line[line_addr][1053] & (~hit)) | (cache_line[k][1053] & (hit));
				cache_line[k][1054] = (mem_line[line_addr][1054] & (~hit)) | (cache_line[k][1054] & (hit));
				cache_line[k][1055] = (mem_line[line_addr][1055] & (~hit)) | (cache_line[k][1055] & (hit));
				cache_line[k][1056] = (mem_line[line_addr][1056] & (~hit)) | (cache_line[k][1056] & (hit));
				cache_line[k][1057] = (mem_line[line_addr][1057] & (~hit)) | (cache_line[k][1057] & (hit));
				cache_line[k][1058] = (mem_line[line_addr][1058] & (~hit)) | (cache_line[k][1058] & (hit));
				cache_line[k][1059] = (mem_line[line_addr][1059] & (~hit)) | (cache_line[k][1059] & (hit));
				cache_line[k][1060] = (mem_line[line_addr][1060] & (~hit)) | (cache_line[k][1060] & (hit));
				cache_line[k][1061] = (mem_line[line_addr][1061] & (~hit)) | (cache_line[k][1061] & (hit));
				cache_line[k][1062] = (mem_line[line_addr][1062] & (~hit)) | (cache_line[k][1062] & (hit));
				cache_line[k][1063] = (mem_line[line_addr][1063] & (~hit)) | (cache_line[k][1063] & (hit));
				cache_line[k][1064] = (mem_line[line_addr][1064] & (~hit)) | (cache_line[k][1064] & (hit));
				cache_line[k][1065] = (mem_line[line_addr][1065] & (~hit)) | (cache_line[k][1065] & (hit));
				cache_line[k][1066] = (mem_line[line_addr][1066] & (~hit)) | (cache_line[k][1066] & (hit));
				cache_line[k][1067] = (mem_line[line_addr][1067] & (~hit)) | (cache_line[k][1067] & (hit));
				cache_line[k][1068] = (mem_line[line_addr][1068] & (~hit)) | (cache_line[k][1068] & (hit));
				cache_line[k][1069] = (mem_line[line_addr][1069] & (~hit)) | (cache_line[k][1069] & (hit));
				cache_line[k][1070] = (mem_line[line_addr][1070] & (~hit)) | (cache_line[k][1070] & (hit));
				cache_line[k][1071] = (mem_line[line_addr][1071] & (~hit)) | (cache_line[k][1071] & (hit));
				cache_line[k][1072] = (mem_line[line_addr][1072] & (~hit)) | (cache_line[k][1072] & (hit));
				cache_line[k][1073] = (mem_line[line_addr][1073] & (~hit)) | (cache_line[k][1073] & (hit));
				cache_line[k][1074] = (mem_line[line_addr][1074] & (~hit)) | (cache_line[k][1074] & (hit));
				cache_line[k][1075] = (mem_line[line_addr][1075] & (~hit)) | (cache_line[k][1075] & (hit));
				cache_line[k][1076] = (mem_line[line_addr][1076] & (~hit)) | (cache_line[k][1076] & (hit));
				cache_line[k][1077] = (mem_line[line_addr][1077] & (~hit)) | (cache_line[k][1077] & (hit));
				cache_line[k][1078] = (mem_line[line_addr][1078] & (~hit)) | (cache_line[k][1078] & (hit));
				cache_line[k][1079] = (mem_line[line_addr][1079] & (~hit)) | (cache_line[k][1079] & (hit));
				cache_line[k][1080] = (mem_line[line_addr][1080] & (~hit)) | (cache_line[k][1080] & (hit));
				cache_line[k][1081] = (mem_line[line_addr][1081] & (~hit)) | (cache_line[k][1081] & (hit));
				cache_line[k][1082] = (mem_line[line_addr][1082] & (~hit)) | (cache_line[k][1082] & (hit));
				cache_line[k][1083] = (mem_line[line_addr][1083] & (~hit)) | (cache_line[k][1083] & (hit));
				cache_line[k][1084] = (mem_line[line_addr][1084] & (~hit)) | (cache_line[k][1084] & (hit));
				cache_line[k][1085] = (mem_line[line_addr][1085] & (~hit)) | (cache_line[k][1085] & (hit));
				cache_line[k][1086] = (mem_line[line_addr][1086] & (~hit)) | (cache_line[k][1086] & (hit));
				cache_line[k][1087] = (mem_line[line_addr][1087] & (~hit)) | (cache_line[k][1087] & (hit));
				cache_line[k][1088] = (mem_line[line_addr][1088] & (~hit)) | (cache_line[k][1088] & (hit));
				cache_line[k][1089] = (mem_line[line_addr][1089] & (~hit)) | (cache_line[k][1089] & (hit));
				cache_line[k][1090] = (mem_line[line_addr][1090] & (~hit)) | (cache_line[k][1090] & (hit));
				cache_line[k][1091] = (mem_line[line_addr][1091] & (~hit)) | (cache_line[k][1091] & (hit));
				cache_line[k][1092] = (mem_line[line_addr][1092] & (~hit)) | (cache_line[k][1092] & (hit));
				cache_line[k][1093] = (mem_line[line_addr][1093] & (~hit)) | (cache_line[k][1093] & (hit));
				cache_line[k][1094] = (mem_line[line_addr][1094] & (~hit)) | (cache_line[k][1094] & (hit));
				cache_line[k][1095] = (mem_line[line_addr][1095] & (~hit)) | (cache_line[k][1095] & (hit));
				cache_line[k][1096] = (mem_line[line_addr][1096] & (~hit)) | (cache_line[k][1096] & (hit));
				cache_line[k][1097] = (mem_line[line_addr][1097] & (~hit)) | (cache_line[k][1097] & (hit));
				cache_line[k][1098] = (mem_line[line_addr][1098] & (~hit)) | (cache_line[k][1098] & (hit));
				cache_line[k][1099] = (mem_line[line_addr][1099] & (~hit)) | (cache_line[k][1099] & (hit));
				cache_line[k][1100] = (mem_line[line_addr][1100] & (~hit)) | (cache_line[k][1100] & (hit));
				cache_line[k][1101] = (mem_line[line_addr][1101] & (~hit)) | (cache_line[k][1101] & (hit));
				cache_line[k][1102] = (mem_line[line_addr][1102] & (~hit)) | (cache_line[k][1102] & (hit));
				cache_line[k][1103] = (mem_line[line_addr][1103] & (~hit)) | (cache_line[k][1103] & (hit));
				cache_line[k][1104] = (mem_line[line_addr][1104] & (~hit)) | (cache_line[k][1104] & (hit));
				cache_line[k][1105] = (mem_line[line_addr][1105] & (~hit)) | (cache_line[k][1105] & (hit));
				cache_line[k][1106] = (mem_line[line_addr][1106] & (~hit)) | (cache_line[k][1106] & (hit));
				cache_line[k][1107] = (mem_line[line_addr][1107] & (~hit)) | (cache_line[k][1107] & (hit));
				cache_line[k][1108] = (mem_line[line_addr][1108] & (~hit)) | (cache_line[k][1108] & (hit));
				cache_line[k][1109] = (mem_line[line_addr][1109] & (~hit)) | (cache_line[k][1109] & (hit));
				cache_line[k][1110] = (mem_line[line_addr][1110] & (~hit)) | (cache_line[k][1110] & (hit));
				cache_line[k][1111] = (mem_line[line_addr][1111] & (~hit)) | (cache_line[k][1111] & (hit));
				cache_line[k][1112] = (mem_line[line_addr][1112] & (~hit)) | (cache_line[k][1112] & (hit));
				cache_line[k][1113] = (mem_line[line_addr][1113] & (~hit)) | (cache_line[k][1113] & (hit));
				cache_line[k][1114] = (mem_line[line_addr][1114] & (~hit)) | (cache_line[k][1114] & (hit));
				cache_line[k][1115] = (mem_line[line_addr][1115] & (~hit)) | (cache_line[k][1115] & (hit));
				cache_line[k][1116] = (mem_line[line_addr][1116] & (~hit)) | (cache_line[k][1116] & (hit));
				cache_line[k][1117] = (mem_line[line_addr][1117] & (~hit)) | (cache_line[k][1117] & (hit));
				cache_line[k][1118] = (mem_line[line_addr][1118] & (~hit)) | (cache_line[k][1118] & (hit));
				cache_line[k][1119] = (mem_line[line_addr][1119] & (~hit)) | (cache_line[k][1119] & (hit));
				cache_line[k][1120] = (mem_line[line_addr][1120] & (~hit)) | (cache_line[k][1120] & (hit));
				cache_line[k][1121] = (mem_line[line_addr][1121] & (~hit)) | (cache_line[k][1121] & (hit));
				cache_line[k][1122] = (mem_line[line_addr][1122] & (~hit)) | (cache_line[k][1122] & (hit));
				cache_line[k][1123] = (mem_line[line_addr][1123] & (~hit)) | (cache_line[k][1123] & (hit));
				cache_line[k][1124] = (mem_line[line_addr][1124] & (~hit)) | (cache_line[k][1124] & (hit));
				cache_line[k][1125] = (mem_line[line_addr][1125] & (~hit)) | (cache_line[k][1125] & (hit));
				cache_line[k][1126] = (mem_line[line_addr][1126] & (~hit)) | (cache_line[k][1126] & (hit));
				cache_line[k][1127] = (mem_line[line_addr][1127] & (~hit)) | (cache_line[k][1127] & (hit));
				cache_line[k][1128] = (mem_line[line_addr][1128] & (~hit)) | (cache_line[k][1128] & (hit));
				cache_line[k][1129] = (mem_line[line_addr][1129] & (~hit)) | (cache_line[k][1129] & (hit));
				cache_line[k][1130] = (mem_line[line_addr][1130] & (~hit)) | (cache_line[k][1130] & (hit));
				cache_line[k][1131] = (mem_line[line_addr][1131] & (~hit)) | (cache_line[k][1131] & (hit));
				cache_line[k][1132] = (mem_line[line_addr][1132] & (~hit)) | (cache_line[k][1132] & (hit));
				cache_line[k][1133] = (mem_line[line_addr][1133] & (~hit)) | (cache_line[k][1133] & (hit));
				cache_line[k][1134] = (mem_line[line_addr][1134] & (~hit)) | (cache_line[k][1134] & (hit));
				cache_line[k][1135] = (mem_line[line_addr][1135] & (~hit)) | (cache_line[k][1135] & (hit));
				cache_line[k][1136] = (mem_line[line_addr][1136] & (~hit)) | (cache_line[k][1136] & (hit));
				cache_line[k][1137] = (mem_line[line_addr][1137] & (~hit)) | (cache_line[k][1137] & (hit));
				cache_line[k][1138] = (mem_line[line_addr][1138] & (~hit)) | (cache_line[k][1138] & (hit));
				cache_line[k][1139] = (mem_line[line_addr][1139] & (~hit)) | (cache_line[k][1139] & (hit));
				cache_line[k][1140] = (mem_line[line_addr][1140] & (~hit)) | (cache_line[k][1140] & (hit));
				cache_line[k][1141] = (mem_line[line_addr][1141] & (~hit)) | (cache_line[k][1141] & (hit));
				cache_line[k][1142] = (mem_line[line_addr][1142] & (~hit)) | (cache_line[k][1142] & (hit));
				cache_line[k][1143] = (mem_line[line_addr][1143] & (~hit)) | (cache_line[k][1143] & (hit));
				cache_line[k][1144] = (mem_line[line_addr][1144] & (~hit)) | (cache_line[k][1144] & (hit));
				cache_line[k][1145] = (mem_line[line_addr][1145] & (~hit)) | (cache_line[k][1145] & (hit));
				cache_line[k][1146] = (mem_line[line_addr][1146] & (~hit)) | (cache_line[k][1146] & (hit));
				cache_line[k][1147] = (mem_line[line_addr][1147] & (~hit)) | (cache_line[k][1147] & (hit));
				cache_line[k][1148] = (mem_line[line_addr][1148] & (~hit)) | (cache_line[k][1148] & (hit));
				cache_line[k][1149] = (mem_line[line_addr][1149] & (~hit)) | (cache_line[k][1149] & (hit));
				cache_line[k][1150] = (mem_line[line_addr][1150] & (~hit)) | (cache_line[k][1150] & (hit));
				cache_line[k][1151] = (mem_line[line_addr][1151] & (~hit)) | (cache_line[k][1151] & (hit));
				cache_line[k][1152] = (mem_line[line_addr][1152] & (~hit)) | (cache_line[k][1152] & (hit));
				cache_line[k][1153] = (mem_line[line_addr][1153] & (~hit)) | (cache_line[k][1153] & (hit));
				cache_line[k][1154] = (mem_line[line_addr][1154] & (~hit)) | (cache_line[k][1154] & (hit));
				cache_line[k][1155] = (mem_line[line_addr][1155] & (~hit)) | (cache_line[k][1155] & (hit));
				cache_line[k][1156] = (mem_line[line_addr][1156] & (~hit)) | (cache_line[k][1156] & (hit));
				cache_line[k][1157] = (mem_line[line_addr][1157] & (~hit)) | (cache_line[k][1157] & (hit));
				cache_line[k][1158] = (mem_line[line_addr][1158] & (~hit)) | (cache_line[k][1158] & (hit));
				cache_line[k][1159] = (mem_line[line_addr][1159] & (~hit)) | (cache_line[k][1159] & (hit));
				cache_line[k][1160] = (mem_line[line_addr][1160] & (~hit)) | (cache_line[k][1160] & (hit));
				cache_line[k][1161] = (mem_line[line_addr][1161] & (~hit)) | (cache_line[k][1161] & (hit));
				cache_line[k][1162] = (mem_line[line_addr][1162] & (~hit)) | (cache_line[k][1162] & (hit));
				cache_line[k][1163] = (mem_line[line_addr][1163] & (~hit)) | (cache_line[k][1163] & (hit));
				cache_line[k][1164] = (mem_line[line_addr][1164] & (~hit)) | (cache_line[k][1164] & (hit));
				cache_line[k][1165] = (mem_line[line_addr][1165] & (~hit)) | (cache_line[k][1165] & (hit));
				cache_line[k][1166] = (mem_line[line_addr][1166] & (~hit)) | (cache_line[k][1166] & (hit));
				cache_line[k][1167] = (mem_line[line_addr][1167] & (~hit)) | (cache_line[k][1167] & (hit));
				cache_line[k][1168] = (mem_line[line_addr][1168] & (~hit)) | (cache_line[k][1168] & (hit));
				cache_line[k][1169] = (mem_line[line_addr][1169] & (~hit)) | (cache_line[k][1169] & (hit));
				cache_line[k][1170] = (mem_line[line_addr][1170] & (~hit)) | (cache_line[k][1170] & (hit));
				cache_line[k][1171] = (mem_line[line_addr][1171] & (~hit)) | (cache_line[k][1171] & (hit));
				cache_line[k][1172] = (mem_line[line_addr][1172] & (~hit)) | (cache_line[k][1172] & (hit));
				cache_line[k][1173] = (mem_line[line_addr][1173] & (~hit)) | (cache_line[k][1173] & (hit));
				cache_line[k][1174] = (mem_line[line_addr][1174] & (~hit)) | (cache_line[k][1174] & (hit));
				cache_line[k][1175] = (mem_line[line_addr][1175] & (~hit)) | (cache_line[k][1175] & (hit));
				cache_line[k][1176] = (mem_line[line_addr][1176] & (~hit)) | (cache_line[k][1176] & (hit));
				cache_line[k][1177] = (mem_line[line_addr][1177] & (~hit)) | (cache_line[k][1177] & (hit));
				cache_line[k][1178] = (mem_line[line_addr][1178] & (~hit)) | (cache_line[k][1178] & (hit));
				cache_line[k][1179] = (mem_line[line_addr][1179] & (~hit)) | (cache_line[k][1179] & (hit));
				cache_line[k][1180] = (mem_line[line_addr][1180] & (~hit)) | (cache_line[k][1180] & (hit));
				cache_line[k][1181] = (mem_line[line_addr][1181] & (~hit)) | (cache_line[k][1181] & (hit));
				cache_line[k][1182] = (mem_line[line_addr][1182] & (~hit)) | (cache_line[k][1182] & (hit));
				cache_line[k][1183] = (mem_line[line_addr][1183] & (~hit)) | (cache_line[k][1183] & (hit));
				cache_line[k][1184] = (mem_line[line_addr][1184] & (~hit)) | (cache_line[k][1184] & (hit));
				cache_line[k][1185] = (mem_line[line_addr][1185] & (~hit)) | (cache_line[k][1185] & (hit));
				cache_line[k][1186] = (mem_line[line_addr][1186] & (~hit)) | (cache_line[k][1186] & (hit));
				cache_line[k][1187] = (mem_line[line_addr][1187] & (~hit)) | (cache_line[k][1187] & (hit));
				cache_line[k][1188] = (mem_line[line_addr][1188] & (~hit)) | (cache_line[k][1188] & (hit));
				cache_line[k][1189] = (mem_line[line_addr][1189] & (~hit)) | (cache_line[k][1189] & (hit));
				cache_line[k][1190] = (mem_line[line_addr][1190] & (~hit)) | (cache_line[k][1190] & (hit));
				cache_line[k][1191] = (mem_line[line_addr][1191] & (~hit)) | (cache_line[k][1191] & (hit));
				cache_line[k][1192] = (mem_line[line_addr][1192] & (~hit)) | (cache_line[k][1192] & (hit));
				cache_line[k][1193] = (mem_line[line_addr][1193] & (~hit)) | (cache_line[k][1193] & (hit));
				cache_line[k][1194] = (mem_line[line_addr][1194] & (~hit)) | (cache_line[k][1194] & (hit));
				cache_line[k][1195] = (mem_line[line_addr][1195] & (~hit)) | (cache_line[k][1195] & (hit));
				cache_line[k][1196] = (mem_line[line_addr][1196] & (~hit)) | (cache_line[k][1196] & (hit));
				cache_line[k][1197] = (mem_line[line_addr][1197] & (~hit)) | (cache_line[k][1197] & (hit));
				cache_line[k][1198] = (mem_line[line_addr][1198] & (~hit)) | (cache_line[k][1198] & (hit));
				cache_line[k][1199] = (mem_line[line_addr][1199] & (~hit)) | (cache_line[k][1199] & (hit));
				cache_line[k][1200] = (mem_line[line_addr][1200] & (~hit)) | (cache_line[k][1200] & (hit));
				cache_line[k][1201] = (mem_line[line_addr][1201] & (~hit)) | (cache_line[k][1201] & (hit));
				cache_line[k][1202] = (mem_line[line_addr][1202] & (~hit)) | (cache_line[k][1202] & (hit));
				cache_line[k][1203] = (mem_line[line_addr][1203] & (~hit)) | (cache_line[k][1203] & (hit));
				cache_line[k][1204] = (mem_line[line_addr][1204] & (~hit)) | (cache_line[k][1204] & (hit));
				cache_line[k][1205] = (mem_line[line_addr][1205] & (~hit)) | (cache_line[k][1205] & (hit));
				cache_line[k][1206] = (mem_line[line_addr][1206] & (~hit)) | (cache_line[k][1206] & (hit));
				cache_line[k][1207] = (mem_line[line_addr][1207] & (~hit)) | (cache_line[k][1207] & (hit));
				cache_line[k][1208] = (mem_line[line_addr][1208] & (~hit)) | (cache_line[k][1208] & (hit));
				cache_line[k][1209] = (mem_line[line_addr][1209] & (~hit)) | (cache_line[k][1209] & (hit));
				cache_line[k][1210] = (mem_line[line_addr][1210] & (~hit)) | (cache_line[k][1210] & (hit));
				cache_line[k][1211] = (mem_line[line_addr][1211] & (~hit)) | (cache_line[k][1211] & (hit));
				cache_line[k][1212] = (mem_line[line_addr][1212] & (~hit)) | (cache_line[k][1212] & (hit));
				cache_line[k][1213] = (mem_line[line_addr][1213] & (~hit)) | (cache_line[k][1213] & (hit));
				cache_line[k][1214] = (mem_line[line_addr][1214] & (~hit)) | (cache_line[k][1214] & (hit));
				cache_line[k][1215] = (mem_line[line_addr][1215] & (~hit)) | (cache_line[k][1215] & (hit));
				cache_line[k][1216] = (mem_line[line_addr][1216] & (~hit)) | (cache_line[k][1216] & (hit));
				cache_line[k][1217] = (mem_line[line_addr][1217] & (~hit)) | (cache_line[k][1217] & (hit));
				cache_line[k][1218] = (mem_line[line_addr][1218] & (~hit)) | (cache_line[k][1218] & (hit));
				cache_line[k][1219] = (mem_line[line_addr][1219] & (~hit)) | (cache_line[k][1219] & (hit));
				cache_line[k][1220] = (mem_line[line_addr][1220] & (~hit)) | (cache_line[k][1220] & (hit));
				cache_line[k][1221] = (mem_line[line_addr][1221] & (~hit)) | (cache_line[k][1221] & (hit));
				cache_line[k][1222] = (mem_line[line_addr][1222] & (~hit)) | (cache_line[k][1222] & (hit));
				cache_line[k][1223] = (mem_line[line_addr][1223] & (~hit)) | (cache_line[k][1223] & (hit));
				cache_line[k][1224] = (mem_line[line_addr][1224] & (~hit)) | (cache_line[k][1224] & (hit));
				cache_line[k][1225] = (mem_line[line_addr][1225] & (~hit)) | (cache_line[k][1225] & (hit));
				cache_line[k][1226] = (mem_line[line_addr][1226] & (~hit)) | (cache_line[k][1226] & (hit));
				cache_line[k][1227] = (mem_line[line_addr][1227] & (~hit)) | (cache_line[k][1227] & (hit));
				cache_line[k][1228] = (mem_line[line_addr][1228] & (~hit)) | (cache_line[k][1228] & (hit));
				cache_line[k][1229] = (mem_line[line_addr][1229] & (~hit)) | (cache_line[k][1229] & (hit));
				cache_line[k][1230] = (mem_line[line_addr][1230] & (~hit)) | (cache_line[k][1230] & (hit));
				cache_line[k][1231] = (mem_line[line_addr][1231] & (~hit)) | (cache_line[k][1231] & (hit));
				cache_line[k][1232] = (mem_line[line_addr][1232] & (~hit)) | (cache_line[k][1232] & (hit));
				cache_line[k][1233] = (mem_line[line_addr][1233] & (~hit)) | (cache_line[k][1233] & (hit));
				cache_line[k][1234] = (mem_line[line_addr][1234] & (~hit)) | (cache_line[k][1234] & (hit));
				cache_line[k][1235] = (mem_line[line_addr][1235] & (~hit)) | (cache_line[k][1235] & (hit));
				cache_line[k][1236] = (mem_line[line_addr][1236] & (~hit)) | (cache_line[k][1236] & (hit));
				cache_line[k][1237] = (mem_line[line_addr][1237] & (~hit)) | (cache_line[k][1237] & (hit));
				cache_line[k][1238] = (mem_line[line_addr][1238] & (~hit)) | (cache_line[k][1238] & (hit));
				cache_line[k][1239] = (mem_line[line_addr][1239] & (~hit)) | (cache_line[k][1239] & (hit));
				cache_line[k][1240] = (mem_line[line_addr][1240] & (~hit)) | (cache_line[k][1240] & (hit));
				cache_line[k][1241] = (mem_line[line_addr][1241] & (~hit)) | (cache_line[k][1241] & (hit));
				cache_line[k][1242] = (mem_line[line_addr][1242] & (~hit)) | (cache_line[k][1242] & (hit));
				cache_line[k][1243] = (mem_line[line_addr][1243] & (~hit)) | (cache_line[k][1243] & (hit));
				cache_line[k][1244] = (mem_line[line_addr][1244] & (~hit)) | (cache_line[k][1244] & (hit));
				cache_line[k][1245] = (mem_line[line_addr][1245] & (~hit)) | (cache_line[k][1245] & (hit));
				cache_line[k][1246] = (mem_line[line_addr][1246] & (~hit)) | (cache_line[k][1246] & (hit));
				cache_line[k][1247] = (mem_line[line_addr][1247] & (~hit)) | (cache_line[k][1247] & (hit));
				cache_line[k][1248] = (mem_line[line_addr][1248] & (~hit)) | (cache_line[k][1248] & (hit));
				cache_line[k][1249] = (mem_line[line_addr][1249] & (~hit)) | (cache_line[k][1249] & (hit));
				cache_line[k][1250] = (mem_line[line_addr][1250] & (~hit)) | (cache_line[k][1250] & (hit));
				cache_line[k][1251] = (mem_line[line_addr][1251] & (~hit)) | (cache_line[k][1251] & (hit));
				cache_line[k][1252] = (mem_line[line_addr][1252] & (~hit)) | (cache_line[k][1252] & (hit));
				cache_line[k][1253] = (mem_line[line_addr][1253] & (~hit)) | (cache_line[k][1253] & (hit));
				cache_line[k][1254] = (mem_line[line_addr][1254] & (~hit)) | (cache_line[k][1254] & (hit));
				cache_line[k][1255] = (mem_line[line_addr][1255] & (~hit)) | (cache_line[k][1255] & (hit));
				cache_line[k][1256] = (mem_line[line_addr][1256] & (~hit)) | (cache_line[k][1256] & (hit));
				cache_line[k][1257] = (mem_line[line_addr][1257] & (~hit)) | (cache_line[k][1257] & (hit));
				cache_line[k][1258] = (mem_line[line_addr][1258] & (~hit)) | (cache_line[k][1258] & (hit));
				cache_line[k][1259] = (mem_line[line_addr][1259] & (~hit)) | (cache_line[k][1259] & (hit));
				cache_line[k][1260] = (mem_line[line_addr][1260] & (~hit)) | (cache_line[k][1260] & (hit));
				cache_line[k][1261] = (mem_line[line_addr][1261] & (~hit)) | (cache_line[k][1261] & (hit));
				cache_line[k][1262] = (mem_line[line_addr][1262] & (~hit)) | (cache_line[k][1262] & (hit));
				cache_line[k][1263] = (mem_line[line_addr][1263] & (~hit)) | (cache_line[k][1263] & (hit));
				cache_line[k][1264] = (mem_line[line_addr][1264] & (~hit)) | (cache_line[k][1264] & (hit));
				cache_line[k][1265] = (mem_line[line_addr][1265] & (~hit)) | (cache_line[k][1265] & (hit));
				cache_line[k][1266] = (mem_line[line_addr][1266] & (~hit)) | (cache_line[k][1266] & (hit));
				cache_line[k][1267] = (mem_line[line_addr][1267] & (~hit)) | (cache_line[k][1267] & (hit));
				cache_line[k][1268] = (mem_line[line_addr][1268] & (~hit)) | (cache_line[k][1268] & (hit));
				cache_line[k][1269] = (mem_line[line_addr][1269] & (~hit)) | (cache_line[k][1269] & (hit));
				cache_line[k][1270] = (mem_line[line_addr][1270] & (~hit)) | (cache_line[k][1270] & (hit));
				cache_line[k][1271] = (mem_line[line_addr][1271] & (~hit)) | (cache_line[k][1271] & (hit));
				cache_line[k][1272] = (mem_line[line_addr][1272] & (~hit)) | (cache_line[k][1272] & (hit));
				cache_line[k][1273] = (mem_line[line_addr][1273] & (~hit)) | (cache_line[k][1273] & (hit));
				cache_line[k][1274] = (mem_line[line_addr][1274] & (~hit)) | (cache_line[k][1274] & (hit));
				cache_line[k][1275] = (mem_line[line_addr][1275] & (~hit)) | (cache_line[k][1275] & (hit));
				cache_line[k][1276] = (mem_line[line_addr][1276] & (~hit)) | (cache_line[k][1276] & (hit));
				cache_line[k][1277] = (mem_line[line_addr][1277] & (~hit)) | (cache_line[k][1277] & (hit));
				cache_line[k][1278] = (mem_line[line_addr][1278] & (~hit)) | (cache_line[k][1278] & (hit));
				cache_line[k][1279] = (mem_line[line_addr][1279] & (~hit)) | (cache_line[k][1279] & (hit));
				cache_line[k][1280] = (mem_line[line_addr][1280] & (~hit)) | (cache_line[k][1280] & (hit));
				cache_line[k][1281] = (mem_line[line_addr][1281] & (~hit)) | (cache_line[k][1281] & (hit));
				cache_line[k][1282] = (mem_line[line_addr][1282] & (~hit)) | (cache_line[k][1282] & (hit));
				cache_line[k][1283] = (mem_line[line_addr][1283] & (~hit)) | (cache_line[k][1283] & (hit));
				cache_line[k][1284] = (mem_line[line_addr][1284] & (~hit)) | (cache_line[k][1284] & (hit));
				cache_line[k][1285] = (mem_line[line_addr][1285] & (~hit)) | (cache_line[k][1285] & (hit));
				cache_line[k][1286] = (mem_line[line_addr][1286] & (~hit)) | (cache_line[k][1286] & (hit));
				cache_line[k][1287] = (mem_line[line_addr][1287] & (~hit)) | (cache_line[k][1287] & (hit));
				cache_line[k][1288] = (mem_line[line_addr][1288] & (~hit)) | (cache_line[k][1288] & (hit));
				cache_line[k][1289] = (mem_line[line_addr][1289] & (~hit)) | (cache_line[k][1289] & (hit));
				cache_line[k][1290] = (mem_line[line_addr][1290] & (~hit)) | (cache_line[k][1290] & (hit));
				cache_line[k][1291] = (mem_line[line_addr][1291] & (~hit)) | (cache_line[k][1291] & (hit));
				cache_line[k][1292] = (mem_line[line_addr][1292] & (~hit)) | (cache_line[k][1292] & (hit));
				cache_line[k][1293] = (mem_line[line_addr][1293] & (~hit)) | (cache_line[k][1293] & (hit));
				cache_line[k][1294] = (mem_line[line_addr][1294] & (~hit)) | (cache_line[k][1294] & (hit));
				cache_line[k][1295] = (mem_line[line_addr][1295] & (~hit)) | (cache_line[k][1295] & (hit));
				cache_line[k][1296] = (mem_line[line_addr][1296] & (~hit)) | (cache_line[k][1296] & (hit));
				cache_line[k][1297] = (mem_line[line_addr][1297] & (~hit)) | (cache_line[k][1297] & (hit));
				cache_line[k][1298] = (mem_line[line_addr][1298] & (~hit)) | (cache_line[k][1298] & (hit));
				cache_line[k][1299] = (mem_line[line_addr][1299] & (~hit)) | (cache_line[k][1299] & (hit));
				cache_line[k][1300] = (mem_line[line_addr][1300] & (~hit)) | (cache_line[k][1300] & (hit));
				cache_line[k][1301] = (mem_line[line_addr][1301] & (~hit)) | (cache_line[k][1301] & (hit));
				cache_line[k][1302] = (mem_line[line_addr][1302] & (~hit)) | (cache_line[k][1302] & (hit));
				cache_line[k][1303] = (mem_line[line_addr][1303] & (~hit)) | (cache_line[k][1303] & (hit));
				cache_line[k][1304] = (mem_line[line_addr][1304] & (~hit)) | (cache_line[k][1304] & (hit));
				cache_line[k][1305] = (mem_line[line_addr][1305] & (~hit)) | (cache_line[k][1305] & (hit));
				cache_line[k][1306] = (mem_line[line_addr][1306] & (~hit)) | (cache_line[k][1306] & (hit));
				cache_line[k][1307] = (mem_line[line_addr][1307] & (~hit)) | (cache_line[k][1307] & (hit));
				cache_line[k][1308] = (mem_line[line_addr][1308] & (~hit)) | (cache_line[k][1308] & (hit));
				cache_line[k][1309] = (mem_line[line_addr][1309] & (~hit)) | (cache_line[k][1309] & (hit));
				cache_line[k][1310] = (mem_line[line_addr][1310] & (~hit)) | (cache_line[k][1310] & (hit));
				cache_line[k][1311] = (mem_line[line_addr][1311] & (~hit)) | (cache_line[k][1311] & (hit));
				cache_line[k][1312] = (mem_line[line_addr][1312] & (~hit)) | (cache_line[k][1312] & (hit));
				cache_line[k][1313] = (mem_line[line_addr][1313] & (~hit)) | (cache_line[k][1313] & (hit));
				cache_line[k][1314] = (mem_line[line_addr][1314] & (~hit)) | (cache_line[k][1314] & (hit));
				cache_line[k][1315] = (mem_line[line_addr][1315] & (~hit)) | (cache_line[k][1315] & (hit));
				cache_line[k][1316] = (mem_line[line_addr][1316] & (~hit)) | (cache_line[k][1316] & (hit));
				cache_line[k][1317] = (mem_line[line_addr][1317] & (~hit)) | (cache_line[k][1317] & (hit));
				cache_line[k][1318] = (mem_line[line_addr][1318] & (~hit)) | (cache_line[k][1318] & (hit));
				cache_line[k][1319] = (mem_line[line_addr][1319] & (~hit)) | (cache_line[k][1319] & (hit));
				cache_line[k][1320] = (mem_line[line_addr][1320] & (~hit)) | (cache_line[k][1320] & (hit));
				cache_line[k][1321] = (mem_line[line_addr][1321] & (~hit)) | (cache_line[k][1321] & (hit));
				cache_line[k][1322] = (mem_line[line_addr][1322] & (~hit)) | (cache_line[k][1322] & (hit));
				cache_line[k][1323] = (mem_line[line_addr][1323] & (~hit)) | (cache_line[k][1323] & (hit));
				cache_line[k][1324] = (mem_line[line_addr][1324] & (~hit)) | (cache_line[k][1324] & (hit));
				cache_line[k][1325] = (mem_line[line_addr][1325] & (~hit)) | (cache_line[k][1325] & (hit));
				cache_line[k][1326] = (mem_line[line_addr][1326] & (~hit)) | (cache_line[k][1326] & (hit));
				cache_line[k][1327] = (mem_line[line_addr][1327] & (~hit)) | (cache_line[k][1327] & (hit));
				cache_line[k][1328] = (mem_line[line_addr][1328] & (~hit)) | (cache_line[k][1328] & (hit));
				cache_line[k][1329] = (mem_line[line_addr][1329] & (~hit)) | (cache_line[k][1329] & (hit));
				cache_line[k][1330] = (mem_line[line_addr][1330] & (~hit)) | (cache_line[k][1330] & (hit));
				cache_line[k][1331] = (mem_line[line_addr][1331] & (~hit)) | (cache_line[k][1331] & (hit));
				cache_line[k][1332] = (mem_line[line_addr][1332] & (~hit)) | (cache_line[k][1332] & (hit));
				cache_line[k][1333] = (mem_line[line_addr][1333] & (~hit)) | (cache_line[k][1333] & (hit));
				cache_line[k][1334] = (mem_line[line_addr][1334] & (~hit)) | (cache_line[k][1334] & (hit));
				cache_line[k][1335] = (mem_line[line_addr][1335] & (~hit)) | (cache_line[k][1335] & (hit));
				cache_line[k][1336] = (mem_line[line_addr][1336] & (~hit)) | (cache_line[k][1336] & (hit));
				cache_line[k][1337] = (mem_line[line_addr][1337] & (~hit)) | (cache_line[k][1337] & (hit));
				cache_line[k][1338] = (mem_line[line_addr][1338] & (~hit)) | (cache_line[k][1338] & (hit));
				cache_line[k][1339] = (mem_line[line_addr][1339] & (~hit)) | (cache_line[k][1339] & (hit));
				cache_line[k][1340] = (mem_line[line_addr][1340] & (~hit)) | (cache_line[k][1340] & (hit));
				cache_line[k][1341] = (mem_line[line_addr][1341] & (~hit)) | (cache_line[k][1341] & (hit));
				cache_line[k][1342] = (mem_line[line_addr][1342] & (~hit)) | (cache_line[k][1342] & (hit));
				cache_line[k][1343] = (mem_line[line_addr][1343] & (~hit)) | (cache_line[k][1343] & (hit));
				cache_line[k][1344] = (mem_line[line_addr][1344] & (~hit)) | (cache_line[k][1344] & (hit));
				cache_line[k][1345] = (mem_line[line_addr][1345] & (~hit)) | (cache_line[k][1345] & (hit));
				cache_line[k][1346] = (mem_line[line_addr][1346] & (~hit)) | (cache_line[k][1346] & (hit));
				cache_line[k][1347] = (mem_line[line_addr][1347] & (~hit)) | (cache_line[k][1347] & (hit));
				cache_line[k][1348] = (mem_line[line_addr][1348] & (~hit)) | (cache_line[k][1348] & (hit));
				cache_line[k][1349] = (mem_line[line_addr][1349] & (~hit)) | (cache_line[k][1349] & (hit));
				cache_line[k][1350] = (mem_line[line_addr][1350] & (~hit)) | (cache_line[k][1350] & (hit));
				cache_line[k][1351] = (mem_line[line_addr][1351] & (~hit)) | (cache_line[k][1351] & (hit));
				cache_line[k][1352] = (mem_line[line_addr][1352] & (~hit)) | (cache_line[k][1352] & (hit));
				cache_line[k][1353] = (mem_line[line_addr][1353] & (~hit)) | (cache_line[k][1353] & (hit));
				cache_line[k][1354] = (mem_line[line_addr][1354] & (~hit)) | (cache_line[k][1354] & (hit));
				cache_line[k][1355] = (mem_line[line_addr][1355] & (~hit)) | (cache_line[k][1355] & (hit));
				cache_line[k][1356] = (mem_line[line_addr][1356] & (~hit)) | (cache_line[k][1356] & (hit));
				cache_line[k][1357] = (mem_line[line_addr][1357] & (~hit)) | (cache_line[k][1357] & (hit));
				cache_line[k][1358] = (mem_line[line_addr][1358] & (~hit)) | (cache_line[k][1358] & (hit));
				cache_line[k][1359] = (mem_line[line_addr][1359] & (~hit)) | (cache_line[k][1359] & (hit));
				cache_line[k][1360] = (mem_line[line_addr][1360] & (~hit)) | (cache_line[k][1360] & (hit));
				cache_line[k][1361] = (mem_line[line_addr][1361] & (~hit)) | (cache_line[k][1361] & (hit));
				cache_line[k][1362] = (mem_line[line_addr][1362] & (~hit)) | (cache_line[k][1362] & (hit));
				cache_line[k][1363] = (mem_line[line_addr][1363] & (~hit)) | (cache_line[k][1363] & (hit));
				cache_line[k][1364] = (mem_line[line_addr][1364] & (~hit)) | (cache_line[k][1364] & (hit));
				cache_line[k][1365] = (mem_line[line_addr][1365] & (~hit)) | (cache_line[k][1365] & (hit));
				cache_line[k][1366] = (mem_line[line_addr][1366] & (~hit)) | (cache_line[k][1366] & (hit));
				cache_line[k][1367] = (mem_line[line_addr][1367] & (~hit)) | (cache_line[k][1367] & (hit));
				cache_line[k][1368] = (mem_line[line_addr][1368] & (~hit)) | (cache_line[k][1368] & (hit));
				cache_line[k][1369] = (mem_line[line_addr][1369] & (~hit)) | (cache_line[k][1369] & (hit));
				cache_line[k][1370] = (mem_line[line_addr][1370] & (~hit)) | (cache_line[k][1370] & (hit));
				cache_line[k][1371] = (mem_line[line_addr][1371] & (~hit)) | (cache_line[k][1371] & (hit));
				cache_line[k][1372] = (mem_line[line_addr][1372] & (~hit)) | (cache_line[k][1372] & (hit));
				cache_line[k][1373] = (mem_line[line_addr][1373] & (~hit)) | (cache_line[k][1373] & (hit));
				cache_line[k][1374] = (mem_line[line_addr][1374] & (~hit)) | (cache_line[k][1374] & (hit));
				cache_line[k][1375] = (mem_line[line_addr][1375] & (~hit)) | (cache_line[k][1375] & (hit));
				cache_line[k][1376] = (mem_line[line_addr][1376] & (~hit)) | (cache_line[k][1376] & (hit));
				cache_line[k][1377] = (mem_line[line_addr][1377] & (~hit)) | (cache_line[k][1377] & (hit));
				cache_line[k][1378] = (mem_line[line_addr][1378] & (~hit)) | (cache_line[k][1378] & (hit));
				cache_line[k][1379] = (mem_line[line_addr][1379] & (~hit)) | (cache_line[k][1379] & (hit));
				cache_line[k][1380] = (mem_line[line_addr][1380] & (~hit)) | (cache_line[k][1380] & (hit));
				cache_line[k][1381] = (mem_line[line_addr][1381] & (~hit)) | (cache_line[k][1381] & (hit));
				cache_line[k][1382] = (mem_line[line_addr][1382] & (~hit)) | (cache_line[k][1382] & (hit));
				cache_line[k][1383] = (mem_line[line_addr][1383] & (~hit)) | (cache_line[k][1383] & (hit));
				cache_line[k][1384] = (mem_line[line_addr][1384] & (~hit)) | (cache_line[k][1384] & (hit));
				cache_line[k][1385] = (mem_line[line_addr][1385] & (~hit)) | (cache_line[k][1385] & (hit));
				cache_line[k][1386] = (mem_line[line_addr][1386] & (~hit)) | (cache_line[k][1386] & (hit));
				cache_line[k][1387] = (mem_line[line_addr][1387] & (~hit)) | (cache_line[k][1387] & (hit));
				cache_line[k][1388] = (mem_line[line_addr][1388] & (~hit)) | (cache_line[k][1388] & (hit));
				cache_line[k][1389] = (mem_line[line_addr][1389] & (~hit)) | (cache_line[k][1389] & (hit));
				cache_line[k][1390] = (mem_line[line_addr][1390] & (~hit)) | (cache_line[k][1390] & (hit));
				cache_line[k][1391] = (mem_line[line_addr][1391] & (~hit)) | (cache_line[k][1391] & (hit));
				cache_line[k][1392] = (mem_line[line_addr][1392] & (~hit)) | (cache_line[k][1392] & (hit));
				cache_line[k][1393] = (mem_line[line_addr][1393] & (~hit)) | (cache_line[k][1393] & (hit));
				cache_line[k][1394] = (mem_line[line_addr][1394] & (~hit)) | (cache_line[k][1394] & (hit));
				cache_line[k][1395] = (mem_line[line_addr][1395] & (~hit)) | (cache_line[k][1395] & (hit));
				cache_line[k][1396] = (mem_line[line_addr][1396] & (~hit)) | (cache_line[k][1396] & (hit));
				cache_line[k][1397] = (mem_line[line_addr][1397] & (~hit)) | (cache_line[k][1397] & (hit));
				cache_line[k][1398] = (mem_line[line_addr][1398] & (~hit)) | (cache_line[k][1398] & (hit));
				cache_line[k][1399] = (mem_line[line_addr][1399] & (~hit)) | (cache_line[k][1399] & (hit));
				cache_line[k][1400] = (mem_line[line_addr][1400] & (~hit)) | (cache_line[k][1400] & (hit));
				cache_line[k][1401] = (mem_line[line_addr][1401] & (~hit)) | (cache_line[k][1401] & (hit));
				cache_line[k][1402] = (mem_line[line_addr][1402] & (~hit)) | (cache_line[k][1402] & (hit));
				cache_line[k][1403] = (mem_line[line_addr][1403] & (~hit)) | (cache_line[k][1403] & (hit));
				cache_line[k][1404] = (mem_line[line_addr][1404] & (~hit)) | (cache_line[k][1404] & (hit));
				cache_line[k][1405] = (mem_line[line_addr][1405] & (~hit)) | (cache_line[k][1405] & (hit));
				cache_line[k][1406] = (mem_line[line_addr][1406] & (~hit)) | (cache_line[k][1406] & (hit));
				cache_line[k][1407] = (mem_line[line_addr][1407] & (~hit)) | (cache_line[k][1407] & (hit));
				cache_line[k][1408] = (mem_line[line_addr][1408] & (~hit)) | (cache_line[k][1408] & (hit));
				cache_line[k][1409] = (mem_line[line_addr][1409] & (~hit)) | (cache_line[k][1409] & (hit));
				cache_line[k][1410] = (mem_line[line_addr][1410] & (~hit)) | (cache_line[k][1410] & (hit));
				cache_line[k][1411] = (mem_line[line_addr][1411] & (~hit)) | (cache_line[k][1411] & (hit));
				cache_line[k][1412] = (mem_line[line_addr][1412] & (~hit)) | (cache_line[k][1412] & (hit));
				cache_line[k][1413] = (mem_line[line_addr][1413] & (~hit)) | (cache_line[k][1413] & (hit));
				cache_line[k][1414] = (mem_line[line_addr][1414] & (~hit)) | (cache_line[k][1414] & (hit));
				cache_line[k][1415] = (mem_line[line_addr][1415] & (~hit)) | (cache_line[k][1415] & (hit));
				cache_line[k][1416] = (mem_line[line_addr][1416] & (~hit)) | (cache_line[k][1416] & (hit));
				cache_line[k][1417] = (mem_line[line_addr][1417] & (~hit)) | (cache_line[k][1417] & (hit));
				cache_line[k][1418] = (mem_line[line_addr][1418] & (~hit)) | (cache_line[k][1418] & (hit));
				cache_line[k][1419] = (mem_line[line_addr][1419] & (~hit)) | (cache_line[k][1419] & (hit));
				cache_line[k][1420] = (mem_line[line_addr][1420] & (~hit)) | (cache_line[k][1420] & (hit));
				cache_line[k][1421] = (mem_line[line_addr][1421] & (~hit)) | (cache_line[k][1421] & (hit));
				cache_line[k][1422] = (mem_line[line_addr][1422] & (~hit)) | (cache_line[k][1422] & (hit));
				cache_line[k][1423] = (mem_line[line_addr][1423] & (~hit)) | (cache_line[k][1423] & (hit));
				cache_line[k][1424] = (mem_line[line_addr][1424] & (~hit)) | (cache_line[k][1424] & (hit));
				cache_line[k][1425] = (mem_line[line_addr][1425] & (~hit)) | (cache_line[k][1425] & (hit));
				cache_line[k][1426] = (mem_line[line_addr][1426] & (~hit)) | (cache_line[k][1426] & (hit));
				cache_line[k][1427] = (mem_line[line_addr][1427] & (~hit)) | (cache_line[k][1427] & (hit));
				cache_line[k][1428] = (mem_line[line_addr][1428] & (~hit)) | (cache_line[k][1428] & (hit));
				cache_line[k][1429] = (mem_line[line_addr][1429] & (~hit)) | (cache_line[k][1429] & (hit));
				cache_line[k][1430] = (mem_line[line_addr][1430] & (~hit)) | (cache_line[k][1430] & (hit));
				cache_line[k][1431] = (mem_line[line_addr][1431] & (~hit)) | (cache_line[k][1431] & (hit));
				cache_line[k][1432] = (mem_line[line_addr][1432] & (~hit)) | (cache_line[k][1432] & (hit));
				cache_line[k][1433] = (mem_line[line_addr][1433] & (~hit)) | (cache_line[k][1433] & (hit));
				cache_line[k][1434] = (mem_line[line_addr][1434] & (~hit)) | (cache_line[k][1434] & (hit));
				cache_line[k][1435] = (mem_line[line_addr][1435] & (~hit)) | (cache_line[k][1435] & (hit));
				cache_line[k][1436] = (mem_line[line_addr][1436] & (~hit)) | (cache_line[k][1436] & (hit));
				cache_line[k][1437] = (mem_line[line_addr][1437] & (~hit)) | (cache_line[k][1437] & (hit));
				cache_line[k][1438] = (mem_line[line_addr][1438] & (~hit)) | (cache_line[k][1438] & (hit));
				cache_line[k][1439] = (mem_line[line_addr][1439] & (~hit)) | (cache_line[k][1439] & (hit));
				cache_line[k][1440] = (mem_line[line_addr][1440] & (~hit)) | (cache_line[k][1440] & (hit));
				cache_line[k][1441] = (mem_line[line_addr][1441] & (~hit)) | (cache_line[k][1441] & (hit));
				cache_line[k][1442] = (mem_line[line_addr][1442] & (~hit)) | (cache_line[k][1442] & (hit));
				cache_line[k][1443] = (mem_line[line_addr][1443] & (~hit)) | (cache_line[k][1443] & (hit));
				cache_line[k][1444] = (mem_line[line_addr][1444] & (~hit)) | (cache_line[k][1444] & (hit));
				cache_line[k][1445] = (mem_line[line_addr][1445] & (~hit)) | (cache_line[k][1445] & (hit));
				cache_line[k][1446] = (mem_line[line_addr][1446] & (~hit)) | (cache_line[k][1446] & (hit));
				cache_line[k][1447] = (mem_line[line_addr][1447] & (~hit)) | (cache_line[k][1447] & (hit));
				cache_line[k][1448] = (mem_line[line_addr][1448] & (~hit)) | (cache_line[k][1448] & (hit));
				cache_line[k][1449] = (mem_line[line_addr][1449] & (~hit)) | (cache_line[k][1449] & (hit));
				cache_line[k][1450] = (mem_line[line_addr][1450] & (~hit)) | (cache_line[k][1450] & (hit));
				cache_line[k][1451] = (mem_line[line_addr][1451] & (~hit)) | (cache_line[k][1451] & (hit));
				cache_line[k][1452] = (mem_line[line_addr][1452] & (~hit)) | (cache_line[k][1452] & (hit));
				cache_line[k][1453] = (mem_line[line_addr][1453] & (~hit)) | (cache_line[k][1453] & (hit));
				cache_line[k][1454] = (mem_line[line_addr][1454] & (~hit)) | (cache_line[k][1454] & (hit));
				cache_line[k][1455] = (mem_line[line_addr][1455] & (~hit)) | (cache_line[k][1455] & (hit));
				cache_line[k][1456] = (mem_line[line_addr][1456] & (~hit)) | (cache_line[k][1456] & (hit));
				cache_line[k][1457] = (mem_line[line_addr][1457] & (~hit)) | (cache_line[k][1457] & (hit));
				cache_line[k][1458] = (mem_line[line_addr][1458] & (~hit)) | (cache_line[k][1458] & (hit));
				cache_line[k][1459] = (mem_line[line_addr][1459] & (~hit)) | (cache_line[k][1459] & (hit));
				cache_line[k][1460] = (mem_line[line_addr][1460] & (~hit)) | (cache_line[k][1460] & (hit));
				cache_line[k][1461] = (mem_line[line_addr][1461] & (~hit)) | (cache_line[k][1461] & (hit));
				cache_line[k][1462] = (mem_line[line_addr][1462] & (~hit)) | (cache_line[k][1462] & (hit));
				cache_line[k][1463] = (mem_line[line_addr][1463] & (~hit)) | (cache_line[k][1463] & (hit));
				cache_line[k][1464] = (mem_line[line_addr][1464] & (~hit)) | (cache_line[k][1464] & (hit));
				cache_line[k][1465] = (mem_line[line_addr][1465] & (~hit)) | (cache_line[k][1465] & (hit));
				cache_line[k][1466] = (mem_line[line_addr][1466] & (~hit)) | (cache_line[k][1466] & (hit));
				cache_line[k][1467] = (mem_line[line_addr][1467] & (~hit)) | (cache_line[k][1467] & (hit));
				cache_line[k][1468] = (mem_line[line_addr][1468] & (~hit)) | (cache_line[k][1468] & (hit));
				cache_line[k][1469] = (mem_line[line_addr][1469] & (~hit)) | (cache_line[k][1469] & (hit));
				cache_line[k][1470] = (mem_line[line_addr][1470] & (~hit)) | (cache_line[k][1470] & (hit));
				cache_line[k][1471] = (mem_line[line_addr][1471] & (~hit)) | (cache_line[k][1471] & (hit));
				cache_line[k][1472] = (mem_line[line_addr][1472] & (~hit)) | (cache_line[k][1472] & (hit));
				cache_line[k][1473] = (mem_line[line_addr][1473] & (~hit)) | (cache_line[k][1473] & (hit));
				cache_line[k][1474] = (mem_line[line_addr][1474] & (~hit)) | (cache_line[k][1474] & (hit));
				cache_line[k][1475] = (mem_line[line_addr][1475] & (~hit)) | (cache_line[k][1475] & (hit));
				cache_line[k][1476] = (mem_line[line_addr][1476] & (~hit)) | (cache_line[k][1476] & (hit));
				cache_line[k][1477] = (mem_line[line_addr][1477] & (~hit)) | (cache_line[k][1477] & (hit));
				cache_line[k][1478] = (mem_line[line_addr][1478] & (~hit)) | (cache_line[k][1478] & (hit));
				cache_line[k][1479] = (mem_line[line_addr][1479] & (~hit)) | (cache_line[k][1479] & (hit));
				cache_line[k][1480] = (mem_line[line_addr][1480] & (~hit)) | (cache_line[k][1480] & (hit));
				cache_line[k][1481] = (mem_line[line_addr][1481] & (~hit)) | (cache_line[k][1481] & (hit));
				cache_line[k][1482] = (mem_line[line_addr][1482] & (~hit)) | (cache_line[k][1482] & (hit));
				cache_line[k][1483] = (mem_line[line_addr][1483] & (~hit)) | (cache_line[k][1483] & (hit));
				cache_line[k][1484] = (mem_line[line_addr][1484] & (~hit)) | (cache_line[k][1484] & (hit));
				cache_line[k][1485] = (mem_line[line_addr][1485] & (~hit)) | (cache_line[k][1485] & (hit));
				cache_line[k][1486] = (mem_line[line_addr][1486] & (~hit)) | (cache_line[k][1486] & (hit));
				cache_line[k][1487] = (mem_line[line_addr][1487] & (~hit)) | (cache_line[k][1487] & (hit));
				cache_line[k][1488] = (mem_line[line_addr][1488] & (~hit)) | (cache_line[k][1488] & (hit));
				cache_line[k][1489] = (mem_line[line_addr][1489] & (~hit)) | (cache_line[k][1489] & (hit));
				cache_line[k][1490] = (mem_line[line_addr][1490] & (~hit)) | (cache_line[k][1490] & (hit));
				cache_line[k][1491] = (mem_line[line_addr][1491] & (~hit)) | (cache_line[k][1491] & (hit));
				cache_line[k][1492] = (mem_line[line_addr][1492] & (~hit)) | (cache_line[k][1492] & (hit));
				cache_line[k][1493] = (mem_line[line_addr][1493] & (~hit)) | (cache_line[k][1493] & (hit));
				cache_line[k][1494] = (mem_line[line_addr][1494] & (~hit)) | (cache_line[k][1494] & (hit));
				cache_line[k][1495] = (mem_line[line_addr][1495] & (~hit)) | (cache_line[k][1495] & (hit));
				cache_line[k][1496] = (mem_line[line_addr][1496] & (~hit)) | (cache_line[k][1496] & (hit));
				cache_line[k][1497] = (mem_line[line_addr][1497] & (~hit)) | (cache_line[k][1497] & (hit));
				cache_line[k][1498] = (mem_line[line_addr][1498] & (~hit)) | (cache_line[k][1498] & (hit));
				cache_line[k][1499] = (mem_line[line_addr][1499] & (~hit)) | (cache_line[k][1499] & (hit));
				cache_line[k][1500] = (mem_line[line_addr][1500] & (~hit)) | (cache_line[k][1500] & (hit));
				cache_line[k][1501] = (mem_line[line_addr][1501] & (~hit)) | (cache_line[k][1501] & (hit));
				cache_line[k][1502] = (mem_line[line_addr][1502] & (~hit)) | (cache_line[k][1502] & (hit));
				cache_line[k][1503] = (mem_line[line_addr][1503] & (~hit)) | (cache_line[k][1503] & (hit));
				cache_line[k][1504] = (mem_line[line_addr][1504] & (~hit)) | (cache_line[k][1504] & (hit));
				cache_line[k][1505] = (mem_line[line_addr][1505] & (~hit)) | (cache_line[k][1505] & (hit));
				cache_line[k][1506] = (mem_line[line_addr][1506] & (~hit)) | (cache_line[k][1506] & (hit));
				cache_line[k][1507] = (mem_line[line_addr][1507] & (~hit)) | (cache_line[k][1507] & (hit));
				cache_line[k][1508] = (mem_line[line_addr][1508] & (~hit)) | (cache_line[k][1508] & (hit));
				cache_line[k][1509] = (mem_line[line_addr][1509] & (~hit)) | (cache_line[k][1509] & (hit));
				cache_line[k][1510] = (mem_line[line_addr][1510] & (~hit)) | (cache_line[k][1510] & (hit));
				cache_line[k][1511] = (mem_line[line_addr][1511] & (~hit)) | (cache_line[k][1511] & (hit));
				cache_line[k][1512] = (mem_line[line_addr][1512] & (~hit)) | (cache_line[k][1512] & (hit));
				cache_line[k][1513] = (mem_line[line_addr][1513] & (~hit)) | (cache_line[k][1513] & (hit));
				cache_line[k][1514] = (mem_line[line_addr][1514] & (~hit)) | (cache_line[k][1514] & (hit));
				cache_line[k][1515] = (mem_line[line_addr][1515] & (~hit)) | (cache_line[k][1515] & (hit));
				cache_line[k][1516] = (mem_line[line_addr][1516] & (~hit)) | (cache_line[k][1516] & (hit));
				cache_line[k][1517] = (mem_line[line_addr][1517] & (~hit)) | (cache_line[k][1517] & (hit));
				cache_line[k][1518] = (mem_line[line_addr][1518] & (~hit)) | (cache_line[k][1518] & (hit));
				cache_line[k][1519] = (mem_line[line_addr][1519] & (~hit)) | (cache_line[k][1519] & (hit));
				cache_line[k][1520] = (mem_line[line_addr][1520] & (~hit)) | (cache_line[k][1520] & (hit));
				cache_line[k][1521] = (mem_line[line_addr][1521] & (~hit)) | (cache_line[k][1521] & (hit));
				cache_line[k][1522] = (mem_line[line_addr][1522] & (~hit)) | (cache_line[k][1522] & (hit));
				cache_line[k][1523] = (mem_line[line_addr][1523] & (~hit)) | (cache_line[k][1523] & (hit));
				cache_line[k][1524] = (mem_line[line_addr][1524] & (~hit)) | (cache_line[k][1524] & (hit));
				cache_line[k][1525] = (mem_line[line_addr][1525] & (~hit)) | (cache_line[k][1525] & (hit));
				cache_line[k][1526] = (mem_line[line_addr][1526] & (~hit)) | (cache_line[k][1526] & (hit));
				cache_line[k][1527] = (mem_line[line_addr][1527] & (~hit)) | (cache_line[k][1527] & (hit));
				cache_line[k][1528] = (mem_line[line_addr][1528] & (~hit)) | (cache_line[k][1528] & (hit));
				cache_line[k][1529] = (mem_line[line_addr][1529] & (~hit)) | (cache_line[k][1529] & (hit));
				cache_line[k][1530] = (mem_line[line_addr][1530] & (~hit)) | (cache_line[k][1530] & (hit));
				cache_line[k][1531] = (mem_line[line_addr][1531] & (~hit)) | (cache_line[k][1531] & (hit));
				cache_line[k][1532] = (mem_line[line_addr][1532] & (~hit)) | (cache_line[k][1532] & (hit));
				cache_line[k][1533] = (mem_line[line_addr][1533] & (~hit)) | (cache_line[k][1533] & (hit));
				cache_line[k][1534] = (mem_line[line_addr][1534] & (~hit)) | (cache_line[k][1534] & (hit));
				cache_line[k][1535] = (mem_line[line_addr][1535] & (~hit)) | (cache_line[k][1535] & (hit));
				cache_line[k][1536] = (mem_line[line_addr][1536] & (~hit)) | (cache_line[k][1536] & (hit));
				cache_line[k][1537] = (mem_line[line_addr][1537] & (~hit)) | (cache_line[k][1537] & (hit));
				cache_line[k][1538] = (mem_line[line_addr][1538] & (~hit)) | (cache_line[k][1538] & (hit));
				cache_line[k][1539] = (mem_line[line_addr][1539] & (~hit)) | (cache_line[k][1539] & (hit));
				cache_line[k][1540] = (mem_line[line_addr][1540] & (~hit)) | (cache_line[k][1540] & (hit));
				cache_line[k][1541] = (mem_line[line_addr][1541] & (~hit)) | (cache_line[k][1541] & (hit));
				cache_line[k][1542] = (mem_line[line_addr][1542] & (~hit)) | (cache_line[k][1542] & (hit));
				cache_line[k][1543] = (mem_line[line_addr][1543] & (~hit)) | (cache_line[k][1543] & (hit));
				cache_line[k][1544] = (mem_line[line_addr][1544] & (~hit)) | (cache_line[k][1544] & (hit));
				cache_line[k][1545] = (mem_line[line_addr][1545] & (~hit)) | (cache_line[k][1545] & (hit));
				cache_line[k][1546] = (mem_line[line_addr][1546] & (~hit)) | (cache_line[k][1546] & (hit));
				cache_line[k][1547] = (mem_line[line_addr][1547] & (~hit)) | (cache_line[k][1547] & (hit));
				cache_line[k][1548] = (mem_line[line_addr][1548] & (~hit)) | (cache_line[k][1548] & (hit));
				cache_line[k][1549] = (mem_line[line_addr][1549] & (~hit)) | (cache_line[k][1549] & (hit));
				cache_line[k][1550] = (mem_line[line_addr][1550] & (~hit)) | (cache_line[k][1550] & (hit));
				cache_line[k][1551] = (mem_line[line_addr][1551] & (~hit)) | (cache_line[k][1551] & (hit));
				cache_line[k][1552] = (mem_line[line_addr][1552] & (~hit)) | (cache_line[k][1552] & (hit));
				cache_line[k][1553] = (mem_line[line_addr][1553] & (~hit)) | (cache_line[k][1553] & (hit));
				cache_line[k][1554] = (mem_line[line_addr][1554] & (~hit)) | (cache_line[k][1554] & (hit));
				cache_line[k][1555] = (mem_line[line_addr][1555] & (~hit)) | (cache_line[k][1555] & (hit));
				cache_line[k][1556] = (mem_line[line_addr][1556] & (~hit)) | (cache_line[k][1556] & (hit));
				cache_line[k][1557] = (mem_line[line_addr][1557] & (~hit)) | (cache_line[k][1557] & (hit));
				cache_line[k][1558] = (mem_line[line_addr][1558] & (~hit)) | (cache_line[k][1558] & (hit));
				cache_line[k][1559] = (mem_line[line_addr][1559] & (~hit)) | (cache_line[k][1559] & (hit));
				cache_line[k][1560] = (mem_line[line_addr][1560] & (~hit)) | (cache_line[k][1560] & (hit));
				cache_line[k][1561] = (mem_line[line_addr][1561] & (~hit)) | (cache_line[k][1561] & (hit));
				cache_line[k][1562] = (mem_line[line_addr][1562] & (~hit)) | (cache_line[k][1562] & (hit));
				cache_line[k][1563] = (mem_line[line_addr][1563] & (~hit)) | (cache_line[k][1563] & (hit));
				cache_line[k][1564] = (mem_line[line_addr][1564] & (~hit)) | (cache_line[k][1564] & (hit));
				cache_line[k][1565] = (mem_line[line_addr][1565] & (~hit)) | (cache_line[k][1565] & (hit));
				cache_line[k][1566] = (mem_line[line_addr][1566] & (~hit)) | (cache_line[k][1566] & (hit));
				cache_line[k][1567] = (mem_line[line_addr][1567] & (~hit)) | (cache_line[k][1567] & (hit));
				cache_line[k][1568] = (mem_line[line_addr][1568] & (~hit)) | (cache_line[k][1568] & (hit));
				cache_line[k][1569] = (mem_line[line_addr][1569] & (~hit)) | (cache_line[k][1569] & (hit));
				cache_line[k][1570] = (mem_line[line_addr][1570] & (~hit)) | (cache_line[k][1570] & (hit));
				cache_line[k][1571] = (mem_line[line_addr][1571] & (~hit)) | (cache_line[k][1571] & (hit));
				cache_line[k][1572] = (mem_line[line_addr][1572] & (~hit)) | (cache_line[k][1572] & (hit));
				cache_line[k][1573] = (mem_line[line_addr][1573] & (~hit)) | (cache_line[k][1573] & (hit));
				cache_line[k][1574] = (mem_line[line_addr][1574] & (~hit)) | (cache_line[k][1574] & (hit));
				cache_line[k][1575] = (mem_line[line_addr][1575] & (~hit)) | (cache_line[k][1575] & (hit));
				cache_line[k][1576] = (mem_line[line_addr][1576] & (~hit)) | (cache_line[k][1576] & (hit));
				cache_line[k][1577] = (mem_line[line_addr][1577] & (~hit)) | (cache_line[k][1577] & (hit));
				cache_line[k][1578] = (mem_line[line_addr][1578] & (~hit)) | (cache_line[k][1578] & (hit));
				cache_line[k][1579] = (mem_line[line_addr][1579] & (~hit)) | (cache_line[k][1579] & (hit));
				cache_line[k][1580] = (mem_line[line_addr][1580] & (~hit)) | (cache_line[k][1580] & (hit));
				cache_line[k][1581] = (mem_line[line_addr][1581] & (~hit)) | (cache_line[k][1581] & (hit));
				cache_line[k][1582] = (mem_line[line_addr][1582] & (~hit)) | (cache_line[k][1582] & (hit));
				cache_line[k][1583] = (mem_line[line_addr][1583] & (~hit)) | (cache_line[k][1583] & (hit));
				cache_line[k][1584] = (mem_line[line_addr][1584] & (~hit)) | (cache_line[k][1584] & (hit));
				cache_line[k][1585] = (mem_line[line_addr][1585] & (~hit)) | (cache_line[k][1585] & (hit));
				cache_line[k][1586] = (mem_line[line_addr][1586] & (~hit)) | (cache_line[k][1586] & (hit));
				cache_line[k][1587] = (mem_line[line_addr][1587] & (~hit)) | (cache_line[k][1587] & (hit));
				cache_line[k][1588] = (mem_line[line_addr][1588] & (~hit)) | (cache_line[k][1588] & (hit));
				cache_line[k][1589] = (mem_line[line_addr][1589] & (~hit)) | (cache_line[k][1589] & (hit));
				cache_line[k][1590] = (mem_line[line_addr][1590] & (~hit)) | (cache_line[k][1590] & (hit));
				cache_line[k][1591] = (mem_line[line_addr][1591] & (~hit)) | (cache_line[k][1591] & (hit));
				cache_line[k][1592] = (mem_line[line_addr][1592] & (~hit)) | (cache_line[k][1592] & (hit));
				cache_line[k][1593] = (mem_line[line_addr][1593] & (~hit)) | (cache_line[k][1593] & (hit));
				cache_line[k][1594] = (mem_line[line_addr][1594] & (~hit)) | (cache_line[k][1594] & (hit));
				cache_line[k][1595] = (mem_line[line_addr][1595] & (~hit)) | (cache_line[k][1595] & (hit));
				cache_line[k][1596] = (mem_line[line_addr][1596] & (~hit)) | (cache_line[k][1596] & (hit));
				cache_line[k][1597] = (mem_line[line_addr][1597] & (~hit)) | (cache_line[k][1597] & (hit));
				cache_line[k][1598] = (mem_line[line_addr][1598] & (~hit)) | (cache_line[k][1598] & (hit));
				cache_line[k][1599] = (mem_line[line_addr][1599] & (~hit)) | (cache_line[k][1599] & (hit));
				cache_line[k][1600] = (mem_line[line_addr][1600] & (~hit)) | (cache_line[k][1600] & (hit));
				cache_line[k][1601] = (mem_line[line_addr][1601] & (~hit)) | (cache_line[k][1601] & (hit));
				cache_line[k][1602] = (mem_line[line_addr][1602] & (~hit)) | (cache_line[k][1602] & (hit));
				cache_line[k][1603] = (mem_line[line_addr][1603] & (~hit)) | (cache_line[k][1603] & (hit));
				cache_line[k][1604] = (mem_line[line_addr][1604] & (~hit)) | (cache_line[k][1604] & (hit));
				cache_line[k][1605] = (mem_line[line_addr][1605] & (~hit)) | (cache_line[k][1605] & (hit));
				cache_line[k][1606] = (mem_line[line_addr][1606] & (~hit)) | (cache_line[k][1606] & (hit));
				cache_line[k][1607] = (mem_line[line_addr][1607] & (~hit)) | (cache_line[k][1607] & (hit));
				cache_line[k][1608] = (mem_line[line_addr][1608] & (~hit)) | (cache_line[k][1608] & (hit));
				cache_line[k][1609] = (mem_line[line_addr][1609] & (~hit)) | (cache_line[k][1609] & (hit));
				cache_line[k][1610] = (mem_line[line_addr][1610] & (~hit)) | (cache_line[k][1610] & (hit));
				cache_line[k][1611] = (mem_line[line_addr][1611] & (~hit)) | (cache_line[k][1611] & (hit));
				cache_line[k][1612] = (mem_line[line_addr][1612] & (~hit)) | (cache_line[k][1612] & (hit));
				cache_line[k][1613] = (mem_line[line_addr][1613] & (~hit)) | (cache_line[k][1613] & (hit));
				cache_line[k][1614] = (mem_line[line_addr][1614] & (~hit)) | (cache_line[k][1614] & (hit));
				cache_line[k][1615] = (mem_line[line_addr][1615] & (~hit)) | (cache_line[k][1615] & (hit));
				cache_line[k][1616] = (mem_line[line_addr][1616] & (~hit)) | (cache_line[k][1616] & (hit));
				cache_line[k][1617] = (mem_line[line_addr][1617] & (~hit)) | (cache_line[k][1617] & (hit));
				cache_line[k][1618] = (mem_line[line_addr][1618] & (~hit)) | (cache_line[k][1618] & (hit));
				cache_line[k][1619] = (mem_line[line_addr][1619] & (~hit)) | (cache_line[k][1619] & (hit));
				cache_line[k][1620] = (mem_line[line_addr][1620] & (~hit)) | (cache_line[k][1620] & (hit));
				cache_line[k][1621] = (mem_line[line_addr][1621] & (~hit)) | (cache_line[k][1621] & (hit));
				cache_line[k][1622] = (mem_line[line_addr][1622] & (~hit)) | (cache_line[k][1622] & (hit));
				cache_line[k][1623] = (mem_line[line_addr][1623] & (~hit)) | (cache_line[k][1623] & (hit));
				cache_line[k][1624] = (mem_line[line_addr][1624] & (~hit)) | (cache_line[k][1624] & (hit));
				cache_line[k][1625] = (mem_line[line_addr][1625] & (~hit)) | (cache_line[k][1625] & (hit));
				cache_line[k][1626] = (mem_line[line_addr][1626] & (~hit)) | (cache_line[k][1626] & (hit));
				cache_line[k][1627] = (mem_line[line_addr][1627] & (~hit)) | (cache_line[k][1627] & (hit));
				cache_line[k][1628] = (mem_line[line_addr][1628] & (~hit)) | (cache_line[k][1628] & (hit));
				cache_line[k][1629] = (mem_line[line_addr][1629] & (~hit)) | (cache_line[k][1629] & (hit));
				cache_line[k][1630] = (mem_line[line_addr][1630] & (~hit)) | (cache_line[k][1630] & (hit));
				cache_line[k][1631] = (mem_line[line_addr][1631] & (~hit)) | (cache_line[k][1631] & (hit));
				cache_line[k][1632] = (mem_line[line_addr][1632] & (~hit)) | (cache_line[k][1632] & (hit));
				cache_line[k][1633] = (mem_line[line_addr][1633] & (~hit)) | (cache_line[k][1633] & (hit));
				cache_line[k][1634] = (mem_line[line_addr][1634] & (~hit)) | (cache_line[k][1634] & (hit));
				cache_line[k][1635] = (mem_line[line_addr][1635] & (~hit)) | (cache_line[k][1635] & (hit));
				cache_line[k][1636] = (mem_line[line_addr][1636] & (~hit)) | (cache_line[k][1636] & (hit));
				cache_line[k][1637] = (mem_line[line_addr][1637] & (~hit)) | (cache_line[k][1637] & (hit));
				cache_line[k][1638] = (mem_line[line_addr][1638] & (~hit)) | (cache_line[k][1638] & (hit));
				cache_line[k][1639] = (mem_line[line_addr][1639] & (~hit)) | (cache_line[k][1639] & (hit));
				cache_line[k][1640] = (mem_line[line_addr][1640] & (~hit)) | (cache_line[k][1640] & (hit));
				cache_line[k][1641] = (mem_line[line_addr][1641] & (~hit)) | (cache_line[k][1641] & (hit));
				cache_line[k][1642] = (mem_line[line_addr][1642] & (~hit)) | (cache_line[k][1642] & (hit));
				cache_line[k][1643] = (mem_line[line_addr][1643] & (~hit)) | (cache_line[k][1643] & (hit));
				cache_line[k][1644] = (mem_line[line_addr][1644] & (~hit)) | (cache_line[k][1644] & (hit));
				cache_line[k][1645] = (mem_line[line_addr][1645] & (~hit)) | (cache_line[k][1645] & (hit));
				cache_line[k][1646] = (mem_line[line_addr][1646] & (~hit)) | (cache_line[k][1646] & (hit));
				cache_line[k][1647] = (mem_line[line_addr][1647] & (~hit)) | (cache_line[k][1647] & (hit));
				cache_line[k][1648] = (mem_line[line_addr][1648] & (~hit)) | (cache_line[k][1648] & (hit));
				cache_line[k][1649] = (mem_line[line_addr][1649] & (~hit)) | (cache_line[k][1649] & (hit));
				cache_line[k][1650] = (mem_line[line_addr][1650] & (~hit)) | (cache_line[k][1650] & (hit));
				cache_line[k][1651] = (mem_line[line_addr][1651] & (~hit)) | (cache_line[k][1651] & (hit));
				cache_line[k][1652] = (mem_line[line_addr][1652] & (~hit)) | (cache_line[k][1652] & (hit));
				cache_line[k][1653] = (mem_line[line_addr][1653] & (~hit)) | (cache_line[k][1653] & (hit));
				cache_line[k][1654] = (mem_line[line_addr][1654] & (~hit)) | (cache_line[k][1654] & (hit));
				cache_line[k][1655] = (mem_line[line_addr][1655] & (~hit)) | (cache_line[k][1655] & (hit));
				cache_line[k][1656] = (mem_line[line_addr][1656] & (~hit)) | (cache_line[k][1656] & (hit));
				cache_line[k][1657] = (mem_line[line_addr][1657] & (~hit)) | (cache_line[k][1657] & (hit));
				cache_line[k][1658] = (mem_line[line_addr][1658] & (~hit)) | (cache_line[k][1658] & (hit));
				cache_line[k][1659] = (mem_line[line_addr][1659] & (~hit)) | (cache_line[k][1659] & (hit));
				cache_line[k][1660] = (mem_line[line_addr][1660] & (~hit)) | (cache_line[k][1660] & (hit));
				cache_line[k][1661] = (mem_line[line_addr][1661] & (~hit)) | (cache_line[k][1661] & (hit));
				cache_line[k][1662] = (mem_line[line_addr][1662] & (~hit)) | (cache_line[k][1662] & (hit));
				cache_line[k][1663] = (mem_line[line_addr][1663] & (~hit)) | (cache_line[k][1663] & (hit));
				cache_line[k][1664] = (mem_line[line_addr][1664] & (~hit)) | (cache_line[k][1664] & (hit));
				cache_line[k][1665] = (mem_line[line_addr][1665] & (~hit)) | (cache_line[k][1665] & (hit));
				cache_line[k][1666] = (mem_line[line_addr][1666] & (~hit)) | (cache_line[k][1666] & (hit));
				cache_line[k][1667] = (mem_line[line_addr][1667] & (~hit)) | (cache_line[k][1667] & (hit));
				cache_line[k][1668] = (mem_line[line_addr][1668] & (~hit)) | (cache_line[k][1668] & (hit));
				cache_line[k][1669] = (mem_line[line_addr][1669] & (~hit)) | (cache_line[k][1669] & (hit));
				cache_line[k][1670] = (mem_line[line_addr][1670] & (~hit)) | (cache_line[k][1670] & (hit));
				cache_line[k][1671] = (mem_line[line_addr][1671] & (~hit)) | (cache_line[k][1671] & (hit));
				cache_line[k][1672] = (mem_line[line_addr][1672] & (~hit)) | (cache_line[k][1672] & (hit));
				cache_line[k][1673] = (mem_line[line_addr][1673] & (~hit)) | (cache_line[k][1673] & (hit));
				cache_line[k][1674] = (mem_line[line_addr][1674] & (~hit)) | (cache_line[k][1674] & (hit));
				cache_line[k][1675] = (mem_line[line_addr][1675] & (~hit)) | (cache_line[k][1675] & (hit));
				cache_line[k][1676] = (mem_line[line_addr][1676] & (~hit)) | (cache_line[k][1676] & (hit));
				cache_line[k][1677] = (mem_line[line_addr][1677] & (~hit)) | (cache_line[k][1677] & (hit));
				cache_line[k][1678] = (mem_line[line_addr][1678] & (~hit)) | (cache_line[k][1678] & (hit));
				cache_line[k][1679] = (mem_line[line_addr][1679] & (~hit)) | (cache_line[k][1679] & (hit));
				cache_line[k][1680] = (mem_line[line_addr][1680] & (~hit)) | (cache_line[k][1680] & (hit));
				cache_line[k][1681] = (mem_line[line_addr][1681] & (~hit)) | (cache_line[k][1681] & (hit));
				cache_line[k][1682] = (mem_line[line_addr][1682] & (~hit)) | (cache_line[k][1682] & (hit));
				cache_line[k][1683] = (mem_line[line_addr][1683] & (~hit)) | (cache_line[k][1683] & (hit));
				cache_line[k][1684] = (mem_line[line_addr][1684] & (~hit)) | (cache_line[k][1684] & (hit));
				cache_line[k][1685] = (mem_line[line_addr][1685] & (~hit)) | (cache_line[k][1685] & (hit));
				cache_line[k][1686] = (mem_line[line_addr][1686] & (~hit)) | (cache_line[k][1686] & (hit));
				cache_line[k][1687] = (mem_line[line_addr][1687] & (~hit)) | (cache_line[k][1687] & (hit));
				cache_line[k][1688] = (mem_line[line_addr][1688] & (~hit)) | (cache_line[k][1688] & (hit));
				cache_line[k][1689] = (mem_line[line_addr][1689] & (~hit)) | (cache_line[k][1689] & (hit));
				cache_line[k][1690] = (mem_line[line_addr][1690] & (~hit)) | (cache_line[k][1690] & (hit));
				cache_line[k][1691] = (mem_line[line_addr][1691] & (~hit)) | (cache_line[k][1691] & (hit));
				cache_line[k][1692] = (mem_line[line_addr][1692] & (~hit)) | (cache_line[k][1692] & (hit));
				cache_line[k][1693] = (mem_line[line_addr][1693] & (~hit)) | (cache_line[k][1693] & (hit));
				cache_line[k][1694] = (mem_line[line_addr][1694] & (~hit)) | (cache_line[k][1694] & (hit));
				cache_line[k][1695] = (mem_line[line_addr][1695] & (~hit)) | (cache_line[k][1695] & (hit));
				cache_line[k][1696] = (mem_line[line_addr][1696] & (~hit)) | (cache_line[k][1696] & (hit));
				cache_line[k][1697] = (mem_line[line_addr][1697] & (~hit)) | (cache_line[k][1697] & (hit));
				cache_line[k][1698] = (mem_line[line_addr][1698] & (~hit)) | (cache_line[k][1698] & (hit));
				cache_line[k][1699] = (mem_line[line_addr][1699] & (~hit)) | (cache_line[k][1699] & (hit));
				cache_line[k][1700] = (mem_line[line_addr][1700] & (~hit)) | (cache_line[k][1700] & (hit));
				cache_line[k][1701] = (mem_line[line_addr][1701] & (~hit)) | (cache_line[k][1701] & (hit));
				cache_line[k][1702] = (mem_line[line_addr][1702] & (~hit)) | (cache_line[k][1702] & (hit));
				cache_line[k][1703] = (mem_line[line_addr][1703] & (~hit)) | (cache_line[k][1703] & (hit));
				cache_line[k][1704] = (mem_line[line_addr][1704] & (~hit)) | (cache_line[k][1704] & (hit));
				cache_line[k][1705] = (mem_line[line_addr][1705] & (~hit)) | (cache_line[k][1705] & (hit));
				cache_line[k][1706] = (mem_line[line_addr][1706] & (~hit)) | (cache_line[k][1706] & (hit));
				cache_line[k][1707] = (mem_line[line_addr][1707] & (~hit)) | (cache_line[k][1707] & (hit));
				cache_line[k][1708] = (mem_line[line_addr][1708] & (~hit)) | (cache_line[k][1708] & (hit));
				cache_line[k][1709] = (mem_line[line_addr][1709] & (~hit)) | (cache_line[k][1709] & (hit));
				cache_line[k][1710] = (mem_line[line_addr][1710] & (~hit)) | (cache_line[k][1710] & (hit));
				cache_line[k][1711] = (mem_line[line_addr][1711] & (~hit)) | (cache_line[k][1711] & (hit));
				cache_line[k][1712] = (mem_line[line_addr][1712] & (~hit)) | (cache_line[k][1712] & (hit));
				cache_line[k][1713] = (mem_line[line_addr][1713] & (~hit)) | (cache_line[k][1713] & (hit));
				cache_line[k][1714] = (mem_line[line_addr][1714] & (~hit)) | (cache_line[k][1714] & (hit));
				cache_line[k][1715] = (mem_line[line_addr][1715] & (~hit)) | (cache_line[k][1715] & (hit));
				cache_line[k][1716] = (mem_line[line_addr][1716] & (~hit)) | (cache_line[k][1716] & (hit));
				cache_line[k][1717] = (mem_line[line_addr][1717] & (~hit)) | (cache_line[k][1717] & (hit));
				cache_line[k][1718] = (mem_line[line_addr][1718] & (~hit)) | (cache_line[k][1718] & (hit));
				cache_line[k][1719] = (mem_line[line_addr][1719] & (~hit)) | (cache_line[k][1719] & (hit));
				cache_line[k][1720] = (mem_line[line_addr][1720] & (~hit)) | (cache_line[k][1720] & (hit));
				cache_line[k][1721] = (mem_line[line_addr][1721] & (~hit)) | (cache_line[k][1721] & (hit));
				cache_line[k][1722] = (mem_line[line_addr][1722] & (~hit)) | (cache_line[k][1722] & (hit));
				cache_line[k][1723] = (mem_line[line_addr][1723] & (~hit)) | (cache_line[k][1723] & (hit));
				cache_line[k][1724] = (mem_line[line_addr][1724] & (~hit)) | (cache_line[k][1724] & (hit));
				cache_line[k][1725] = (mem_line[line_addr][1725] & (~hit)) | (cache_line[k][1725] & (hit));
				cache_line[k][1726] = (mem_line[line_addr][1726] & (~hit)) | (cache_line[k][1726] & (hit));
				cache_line[k][1727] = (mem_line[line_addr][1727] & (~hit)) | (cache_line[k][1727] & (hit));
				cache_line[k][1728] = (mem_line[line_addr][1728] & (~hit)) | (cache_line[k][1728] & (hit));
				cache_line[k][1729] = (mem_line[line_addr][1729] & (~hit)) | (cache_line[k][1729] & (hit));
				cache_line[k][1730] = (mem_line[line_addr][1730] & (~hit)) | (cache_line[k][1730] & (hit));
				cache_line[k][1731] = (mem_line[line_addr][1731] & (~hit)) | (cache_line[k][1731] & (hit));
				cache_line[k][1732] = (mem_line[line_addr][1732] & (~hit)) | (cache_line[k][1732] & (hit));
				cache_line[k][1733] = (mem_line[line_addr][1733] & (~hit)) | (cache_line[k][1733] & (hit));
				cache_line[k][1734] = (mem_line[line_addr][1734] & (~hit)) | (cache_line[k][1734] & (hit));
				cache_line[k][1735] = (mem_line[line_addr][1735] & (~hit)) | (cache_line[k][1735] & (hit));
				cache_line[k][1736] = (mem_line[line_addr][1736] & (~hit)) | (cache_line[k][1736] & (hit));
				cache_line[k][1737] = (mem_line[line_addr][1737] & (~hit)) | (cache_line[k][1737] & (hit));
				cache_line[k][1738] = (mem_line[line_addr][1738] & (~hit)) | (cache_line[k][1738] & (hit));
				cache_line[k][1739] = (mem_line[line_addr][1739] & (~hit)) | (cache_line[k][1739] & (hit));
				cache_line[k][1740] = (mem_line[line_addr][1740] & (~hit)) | (cache_line[k][1740] & (hit));
				cache_line[k][1741] = (mem_line[line_addr][1741] & (~hit)) | (cache_line[k][1741] & (hit));
				cache_line[k][1742] = (mem_line[line_addr][1742] & (~hit)) | (cache_line[k][1742] & (hit));
				cache_line[k][1743] = (mem_line[line_addr][1743] & (~hit)) | (cache_line[k][1743] & (hit));
				cache_line[k][1744] = (mem_line[line_addr][1744] & (~hit)) | (cache_line[k][1744] & (hit));
				cache_line[k][1745] = (mem_line[line_addr][1745] & (~hit)) | (cache_line[k][1745] & (hit));
				cache_line[k][1746] = (mem_line[line_addr][1746] & (~hit)) | (cache_line[k][1746] & (hit));
				cache_line[k][1747] = (mem_line[line_addr][1747] & (~hit)) | (cache_line[k][1747] & (hit));
				cache_line[k][1748] = (mem_line[line_addr][1748] & (~hit)) | (cache_line[k][1748] & (hit));
				cache_line[k][1749] = (mem_line[line_addr][1749] & (~hit)) | (cache_line[k][1749] & (hit));
				cache_line[k][1750] = (mem_line[line_addr][1750] & (~hit)) | (cache_line[k][1750] & (hit));
				cache_line[k][1751] = (mem_line[line_addr][1751] & (~hit)) | (cache_line[k][1751] & (hit));
				cache_line[k][1752] = (mem_line[line_addr][1752] & (~hit)) | (cache_line[k][1752] & (hit));
				cache_line[k][1753] = (mem_line[line_addr][1753] & (~hit)) | (cache_line[k][1753] & (hit));
				cache_line[k][1754] = (mem_line[line_addr][1754] & (~hit)) | (cache_line[k][1754] & (hit));
				cache_line[k][1755] = (mem_line[line_addr][1755] & (~hit)) | (cache_line[k][1755] & (hit));
				cache_line[k][1756] = (mem_line[line_addr][1756] & (~hit)) | (cache_line[k][1756] & (hit));
				cache_line[k][1757] = (mem_line[line_addr][1757] & (~hit)) | (cache_line[k][1757] & (hit));
				cache_line[k][1758] = (mem_line[line_addr][1758] & (~hit)) | (cache_line[k][1758] & (hit));
				cache_line[k][1759] = (mem_line[line_addr][1759] & (~hit)) | (cache_line[k][1759] & (hit));
				cache_line[k][1760] = (mem_line[line_addr][1760] & (~hit)) | (cache_line[k][1760] & (hit));
				cache_line[k][1761] = (mem_line[line_addr][1761] & (~hit)) | (cache_line[k][1761] & (hit));
				cache_line[k][1762] = (mem_line[line_addr][1762] & (~hit)) | (cache_line[k][1762] & (hit));
				cache_line[k][1763] = (mem_line[line_addr][1763] & (~hit)) | (cache_line[k][1763] & (hit));
				cache_line[k][1764] = (mem_line[line_addr][1764] & (~hit)) | (cache_line[k][1764] & (hit));
				cache_line[k][1765] = (mem_line[line_addr][1765] & (~hit)) | (cache_line[k][1765] & (hit));
				cache_line[k][1766] = (mem_line[line_addr][1766] & (~hit)) | (cache_line[k][1766] & (hit));
				cache_line[k][1767] = (mem_line[line_addr][1767] & (~hit)) | (cache_line[k][1767] & (hit));
				cache_line[k][1768] = (mem_line[line_addr][1768] & (~hit)) | (cache_line[k][1768] & (hit));
				cache_line[k][1769] = (mem_line[line_addr][1769] & (~hit)) | (cache_line[k][1769] & (hit));
				cache_line[k][1770] = (mem_line[line_addr][1770] & (~hit)) | (cache_line[k][1770] & (hit));
				cache_line[k][1771] = (mem_line[line_addr][1771] & (~hit)) | (cache_line[k][1771] & (hit));
				cache_line[k][1772] = (mem_line[line_addr][1772] & (~hit)) | (cache_line[k][1772] & (hit));
				cache_line[k][1773] = (mem_line[line_addr][1773] & (~hit)) | (cache_line[k][1773] & (hit));
				cache_line[k][1774] = (mem_line[line_addr][1774] & (~hit)) | (cache_line[k][1774] & (hit));
				cache_line[k][1775] = (mem_line[line_addr][1775] & (~hit)) | (cache_line[k][1775] & (hit));
				cache_line[k][1776] = (mem_line[line_addr][1776] & (~hit)) | (cache_line[k][1776] & (hit));
				cache_line[k][1777] = (mem_line[line_addr][1777] & (~hit)) | (cache_line[k][1777] & (hit));
				cache_line[k][1778] = (mem_line[line_addr][1778] & (~hit)) | (cache_line[k][1778] & (hit));
				cache_line[k][1779] = (mem_line[line_addr][1779] & (~hit)) | (cache_line[k][1779] & (hit));
				cache_line[k][1780] = (mem_line[line_addr][1780] & (~hit)) | (cache_line[k][1780] & (hit));
				cache_line[k][1781] = (mem_line[line_addr][1781] & (~hit)) | (cache_line[k][1781] & (hit));
				cache_line[k][1782] = (mem_line[line_addr][1782] & (~hit)) | (cache_line[k][1782] & (hit));
				cache_line[k][1783] = (mem_line[line_addr][1783] & (~hit)) | (cache_line[k][1783] & (hit));
				cache_line[k][1784] = (mem_line[line_addr][1784] & (~hit)) | (cache_line[k][1784] & (hit));
				cache_line[k][1785] = (mem_line[line_addr][1785] & (~hit)) | (cache_line[k][1785] & (hit));
				cache_line[k][1786] = (mem_line[line_addr][1786] & (~hit)) | (cache_line[k][1786] & (hit));
				cache_line[k][1787] = (mem_line[line_addr][1787] & (~hit)) | (cache_line[k][1787] & (hit));
				cache_line[k][1788] = (mem_line[line_addr][1788] & (~hit)) | (cache_line[k][1788] & (hit));
				cache_line[k][1789] = (mem_line[line_addr][1789] & (~hit)) | (cache_line[k][1789] & (hit));
				cache_line[k][1790] = (mem_line[line_addr][1790] & (~hit)) | (cache_line[k][1790] & (hit));
				cache_line[k][1791] = (mem_line[line_addr][1791] & (~hit)) | (cache_line[k][1791] & (hit));
				cache_line[k][1792] = (mem_line[line_addr][1792] & (~hit)) | (cache_line[k][1792] & (hit));
				cache_line[k][1793] = (mem_line[line_addr][1793] & (~hit)) | (cache_line[k][1793] & (hit));
				cache_line[k][1794] = (mem_line[line_addr][1794] & (~hit)) | (cache_line[k][1794] & (hit));
				cache_line[k][1795] = (mem_line[line_addr][1795] & (~hit)) | (cache_line[k][1795] & (hit));
				cache_line[k][1796] = (mem_line[line_addr][1796] & (~hit)) | (cache_line[k][1796] & (hit));
				cache_line[k][1797] = (mem_line[line_addr][1797] & (~hit)) | (cache_line[k][1797] & (hit));
				cache_line[k][1798] = (mem_line[line_addr][1798] & (~hit)) | (cache_line[k][1798] & (hit));
				cache_line[k][1799] = (mem_line[line_addr][1799] & (~hit)) | (cache_line[k][1799] & (hit));
				cache_line[k][1800] = (mem_line[line_addr][1800] & (~hit)) | (cache_line[k][1800] & (hit));
				cache_line[k][1801] = (mem_line[line_addr][1801] & (~hit)) | (cache_line[k][1801] & (hit));
				cache_line[k][1802] = (mem_line[line_addr][1802] & (~hit)) | (cache_line[k][1802] & (hit));
				cache_line[k][1803] = (mem_line[line_addr][1803] & (~hit)) | (cache_line[k][1803] & (hit));
				cache_line[k][1804] = (mem_line[line_addr][1804] & (~hit)) | (cache_line[k][1804] & (hit));
				cache_line[k][1805] = (mem_line[line_addr][1805] & (~hit)) | (cache_line[k][1805] & (hit));
				cache_line[k][1806] = (mem_line[line_addr][1806] & (~hit)) | (cache_line[k][1806] & (hit));
				cache_line[k][1807] = (mem_line[line_addr][1807] & (~hit)) | (cache_line[k][1807] & (hit));
				cache_line[k][1808] = (mem_line[line_addr][1808] & (~hit)) | (cache_line[k][1808] & (hit));
				cache_line[k][1809] = (mem_line[line_addr][1809] & (~hit)) | (cache_line[k][1809] & (hit));
				cache_line[k][1810] = (mem_line[line_addr][1810] & (~hit)) | (cache_line[k][1810] & (hit));
				cache_line[k][1811] = (mem_line[line_addr][1811] & (~hit)) | (cache_line[k][1811] & (hit));
				cache_line[k][1812] = (mem_line[line_addr][1812] & (~hit)) | (cache_line[k][1812] & (hit));
				cache_line[k][1813] = (mem_line[line_addr][1813] & (~hit)) | (cache_line[k][1813] & (hit));
				cache_line[k][1814] = (mem_line[line_addr][1814] & (~hit)) | (cache_line[k][1814] & (hit));
				cache_line[k][1815] = (mem_line[line_addr][1815] & (~hit)) | (cache_line[k][1815] & (hit));
				cache_line[k][1816] = (mem_line[line_addr][1816] & (~hit)) | (cache_line[k][1816] & (hit));
				cache_line[k][1817] = (mem_line[line_addr][1817] & (~hit)) | (cache_line[k][1817] & (hit));
				cache_line[k][1818] = (mem_line[line_addr][1818] & (~hit)) | (cache_line[k][1818] & (hit));
				cache_line[k][1819] = (mem_line[line_addr][1819] & (~hit)) | (cache_line[k][1819] & (hit));
				cache_line[k][1820] = (mem_line[line_addr][1820] & (~hit)) | (cache_line[k][1820] & (hit));
				cache_line[k][1821] = (mem_line[line_addr][1821] & (~hit)) | (cache_line[k][1821] & (hit));
				cache_line[k][1822] = (mem_line[line_addr][1822] & (~hit)) | (cache_line[k][1822] & (hit));
				cache_line[k][1823] = (mem_line[line_addr][1823] & (~hit)) | (cache_line[k][1823] & (hit));
				cache_line[k][1824] = (mem_line[line_addr][1824] & (~hit)) | (cache_line[k][1824] & (hit));
				cache_line[k][1825] = (mem_line[line_addr][1825] & (~hit)) | (cache_line[k][1825] & (hit));
				cache_line[k][1826] = (mem_line[line_addr][1826] & (~hit)) | (cache_line[k][1826] & (hit));
				cache_line[k][1827] = (mem_line[line_addr][1827] & (~hit)) | (cache_line[k][1827] & (hit));
				cache_line[k][1828] = (mem_line[line_addr][1828] & (~hit)) | (cache_line[k][1828] & (hit));
				cache_line[k][1829] = (mem_line[line_addr][1829] & (~hit)) | (cache_line[k][1829] & (hit));
				cache_line[k][1830] = (mem_line[line_addr][1830] & (~hit)) | (cache_line[k][1830] & (hit));
				cache_line[k][1831] = (mem_line[line_addr][1831] & (~hit)) | (cache_line[k][1831] & (hit));
				cache_line[k][1832] = (mem_line[line_addr][1832] & (~hit)) | (cache_line[k][1832] & (hit));
				cache_line[k][1833] = (mem_line[line_addr][1833] & (~hit)) | (cache_line[k][1833] & (hit));
				cache_line[k][1834] = (mem_line[line_addr][1834] & (~hit)) | (cache_line[k][1834] & (hit));
				cache_line[k][1835] = (mem_line[line_addr][1835] & (~hit)) | (cache_line[k][1835] & (hit));
				cache_line[k][1836] = (mem_line[line_addr][1836] & (~hit)) | (cache_line[k][1836] & (hit));
				cache_line[k][1837] = (mem_line[line_addr][1837] & (~hit)) | (cache_line[k][1837] & (hit));
				cache_line[k][1838] = (mem_line[line_addr][1838] & (~hit)) | (cache_line[k][1838] & (hit));
				cache_line[k][1839] = (mem_line[line_addr][1839] & (~hit)) | (cache_line[k][1839] & (hit));
				cache_line[k][1840] = (mem_line[line_addr][1840] & (~hit)) | (cache_line[k][1840] & (hit));
				cache_line[k][1841] = (mem_line[line_addr][1841] & (~hit)) | (cache_line[k][1841] & (hit));
				cache_line[k][1842] = (mem_line[line_addr][1842] & (~hit)) | (cache_line[k][1842] & (hit));
				cache_line[k][1843] = (mem_line[line_addr][1843] & (~hit)) | (cache_line[k][1843] & (hit));
				cache_line[k][1844] = (mem_line[line_addr][1844] & (~hit)) | (cache_line[k][1844] & (hit));
				cache_line[k][1845] = (mem_line[line_addr][1845] & (~hit)) | (cache_line[k][1845] & (hit));
				cache_line[k][1846] = (mem_line[line_addr][1846] & (~hit)) | (cache_line[k][1846] & (hit));
				cache_line[k][1847] = (mem_line[line_addr][1847] & (~hit)) | (cache_line[k][1847] & (hit));
				cache_line[k][1848] = (mem_line[line_addr][1848] & (~hit)) | (cache_line[k][1848] & (hit));
				cache_line[k][1849] = (mem_line[line_addr][1849] & (~hit)) | (cache_line[k][1849] & (hit));
				cache_line[k][1850] = (mem_line[line_addr][1850] & (~hit)) | (cache_line[k][1850] & (hit));
				cache_line[k][1851] = (mem_line[line_addr][1851] & (~hit)) | (cache_line[k][1851] & (hit));
				cache_line[k][1852] = (mem_line[line_addr][1852] & (~hit)) | (cache_line[k][1852] & (hit));
				cache_line[k][1853] = (mem_line[line_addr][1853] & (~hit)) | (cache_line[k][1853] & (hit));
				cache_line[k][1854] = (mem_line[line_addr][1854] & (~hit)) | (cache_line[k][1854] & (hit));
				cache_line[k][1855] = (mem_line[line_addr][1855] & (~hit)) | (cache_line[k][1855] & (hit));
				cache_line[k][1856] = (mem_line[line_addr][1856] & (~hit)) | (cache_line[k][1856] & (hit));
				cache_line[k][1857] = (mem_line[line_addr][1857] & (~hit)) | (cache_line[k][1857] & (hit));
				cache_line[k][1858] = (mem_line[line_addr][1858] & (~hit)) | (cache_line[k][1858] & (hit));
				cache_line[k][1859] = (mem_line[line_addr][1859] & (~hit)) | (cache_line[k][1859] & (hit));
				cache_line[k][1860] = (mem_line[line_addr][1860] & (~hit)) | (cache_line[k][1860] & (hit));
				cache_line[k][1861] = (mem_line[line_addr][1861] & (~hit)) | (cache_line[k][1861] & (hit));
				cache_line[k][1862] = (mem_line[line_addr][1862] & (~hit)) | (cache_line[k][1862] & (hit));
				cache_line[k][1863] = (mem_line[line_addr][1863] & (~hit)) | (cache_line[k][1863] & (hit));
				cache_line[k][1864] = (mem_line[line_addr][1864] & (~hit)) | (cache_line[k][1864] & (hit));
				cache_line[k][1865] = (mem_line[line_addr][1865] & (~hit)) | (cache_line[k][1865] & (hit));
				cache_line[k][1866] = (mem_line[line_addr][1866] & (~hit)) | (cache_line[k][1866] & (hit));
				cache_line[k][1867] = (mem_line[line_addr][1867] & (~hit)) | (cache_line[k][1867] & (hit));
				cache_line[k][1868] = (mem_line[line_addr][1868] & (~hit)) | (cache_line[k][1868] & (hit));
				cache_line[k][1869] = (mem_line[line_addr][1869] & (~hit)) | (cache_line[k][1869] & (hit));
				cache_line[k][1870] = (mem_line[line_addr][1870] & (~hit)) | (cache_line[k][1870] & (hit));
				cache_line[k][1871] = (mem_line[line_addr][1871] & (~hit)) | (cache_line[k][1871] & (hit));
				cache_line[k][1872] = (mem_line[line_addr][1872] & (~hit)) | (cache_line[k][1872] & (hit));
				cache_line[k][1873] = (mem_line[line_addr][1873] & (~hit)) | (cache_line[k][1873] & (hit));
				cache_line[k][1874] = (mem_line[line_addr][1874] & (~hit)) | (cache_line[k][1874] & (hit));
				cache_line[k][1875] = (mem_line[line_addr][1875] & (~hit)) | (cache_line[k][1875] & (hit));
				cache_line[k][1876] = (mem_line[line_addr][1876] & (~hit)) | (cache_line[k][1876] & (hit));
				cache_line[k][1877] = (mem_line[line_addr][1877] & (~hit)) | (cache_line[k][1877] & (hit));
				cache_line[k][1878] = (mem_line[line_addr][1878] & (~hit)) | (cache_line[k][1878] & (hit));
				cache_line[k][1879] = (mem_line[line_addr][1879] & (~hit)) | (cache_line[k][1879] & (hit));
				cache_line[k][1880] = (mem_line[line_addr][1880] & (~hit)) | (cache_line[k][1880] & (hit));
				cache_line[k][1881] = (mem_line[line_addr][1881] & (~hit)) | (cache_line[k][1881] & (hit));
				cache_line[k][1882] = (mem_line[line_addr][1882] & (~hit)) | (cache_line[k][1882] & (hit));
				cache_line[k][1883] = (mem_line[line_addr][1883] & (~hit)) | (cache_line[k][1883] & (hit));
				cache_line[k][1884] = (mem_line[line_addr][1884] & (~hit)) | (cache_line[k][1884] & (hit));
				cache_line[k][1885] = (mem_line[line_addr][1885] & (~hit)) | (cache_line[k][1885] & (hit));
				cache_line[k][1886] = (mem_line[line_addr][1886] & (~hit)) | (cache_line[k][1886] & (hit));
				cache_line[k][1887] = (mem_line[line_addr][1887] & (~hit)) | (cache_line[k][1887] & (hit));
				cache_line[k][1888] = (mem_line[line_addr][1888] & (~hit)) | (cache_line[k][1888] & (hit));
				cache_line[k][1889] = (mem_line[line_addr][1889] & (~hit)) | (cache_line[k][1889] & (hit));
				cache_line[k][1890] = (mem_line[line_addr][1890] & (~hit)) | (cache_line[k][1890] & (hit));
				cache_line[k][1891] = (mem_line[line_addr][1891] & (~hit)) | (cache_line[k][1891] & (hit));
				cache_line[k][1892] = (mem_line[line_addr][1892] & (~hit)) | (cache_line[k][1892] & (hit));
				cache_line[k][1893] = (mem_line[line_addr][1893] & (~hit)) | (cache_line[k][1893] & (hit));
				cache_line[k][1894] = (mem_line[line_addr][1894] & (~hit)) | (cache_line[k][1894] & (hit));
				cache_line[k][1895] = (mem_line[line_addr][1895] & (~hit)) | (cache_line[k][1895] & (hit));
				cache_line[k][1896] = (mem_line[line_addr][1896] & (~hit)) | (cache_line[k][1896] & (hit));
				cache_line[k][1897] = (mem_line[line_addr][1897] & (~hit)) | (cache_line[k][1897] & (hit));
				cache_line[k][1898] = (mem_line[line_addr][1898] & (~hit)) | (cache_line[k][1898] & (hit));
				cache_line[k][1899] = (mem_line[line_addr][1899] & (~hit)) | (cache_line[k][1899] & (hit));
				cache_line[k][1900] = (mem_line[line_addr][1900] & (~hit)) | (cache_line[k][1900] & (hit));
				cache_line[k][1901] = (mem_line[line_addr][1901] & (~hit)) | (cache_line[k][1901] & (hit));
				cache_line[k][1902] = (mem_line[line_addr][1902] & (~hit)) | (cache_line[k][1902] & (hit));
				cache_line[k][1903] = (mem_line[line_addr][1903] & (~hit)) | (cache_line[k][1903] & (hit));
				cache_line[k][1904] = (mem_line[line_addr][1904] & (~hit)) | (cache_line[k][1904] & (hit));
				cache_line[k][1905] = (mem_line[line_addr][1905] & (~hit)) | (cache_line[k][1905] & (hit));
				cache_line[k][1906] = (mem_line[line_addr][1906] & (~hit)) | (cache_line[k][1906] & (hit));
				cache_line[k][1907] = (mem_line[line_addr][1907] & (~hit)) | (cache_line[k][1907] & (hit));
				cache_line[k][1908] = (mem_line[line_addr][1908] & (~hit)) | (cache_line[k][1908] & (hit));
				cache_line[k][1909] = (mem_line[line_addr][1909] & (~hit)) | (cache_line[k][1909] & (hit));
				cache_line[k][1910] = (mem_line[line_addr][1910] & (~hit)) | (cache_line[k][1910] & (hit));
				cache_line[k][1911] = (mem_line[line_addr][1911] & (~hit)) | (cache_line[k][1911] & (hit));
				cache_line[k][1912] = (mem_line[line_addr][1912] & (~hit)) | (cache_line[k][1912] & (hit));
				cache_line[k][1913] = (mem_line[line_addr][1913] & (~hit)) | (cache_line[k][1913] & (hit));
				cache_line[k][1914] = (mem_line[line_addr][1914] & (~hit)) | (cache_line[k][1914] & (hit));
				cache_line[k][1915] = (mem_line[line_addr][1915] & (~hit)) | (cache_line[k][1915] & (hit));
				cache_line[k][1916] = (mem_line[line_addr][1916] & (~hit)) | (cache_line[k][1916] & (hit));
				cache_line[k][1917] = (mem_line[line_addr][1917] & (~hit)) | (cache_line[k][1917] & (hit));
				cache_line[k][1918] = (mem_line[line_addr][1918] & (~hit)) | (cache_line[k][1918] & (hit));
				cache_line[k][1919] = (mem_line[line_addr][1919] & (~hit)) | (cache_line[k][1919] & (hit));
				cache_line[k][1920] = (mem_line[line_addr][1920] & (~hit)) | (cache_line[k][1920] & (hit));
				cache_line[k][1921] = (mem_line[line_addr][1921] & (~hit)) | (cache_line[k][1921] & (hit));
				cache_line[k][1922] = (mem_line[line_addr][1922] & (~hit)) | (cache_line[k][1922] & (hit));
				cache_line[k][1923] = (mem_line[line_addr][1923] & (~hit)) | (cache_line[k][1923] & (hit));
				cache_line[k][1924] = (mem_line[line_addr][1924] & (~hit)) | (cache_line[k][1924] & (hit));
				cache_line[k][1925] = (mem_line[line_addr][1925] & (~hit)) | (cache_line[k][1925] & (hit));
				cache_line[k][1926] = (mem_line[line_addr][1926] & (~hit)) | (cache_line[k][1926] & (hit));
				cache_line[k][1927] = (mem_line[line_addr][1927] & (~hit)) | (cache_line[k][1927] & (hit));
				cache_line[k][1928] = (mem_line[line_addr][1928] & (~hit)) | (cache_line[k][1928] & (hit));
				cache_line[k][1929] = (mem_line[line_addr][1929] & (~hit)) | (cache_line[k][1929] & (hit));
				cache_line[k][1930] = (mem_line[line_addr][1930] & (~hit)) | (cache_line[k][1930] & (hit));
				cache_line[k][1931] = (mem_line[line_addr][1931] & (~hit)) | (cache_line[k][1931] & (hit));
				cache_line[k][1932] = (mem_line[line_addr][1932] & (~hit)) | (cache_line[k][1932] & (hit));
				cache_line[k][1933] = (mem_line[line_addr][1933] & (~hit)) | (cache_line[k][1933] & (hit));
				cache_line[k][1934] = (mem_line[line_addr][1934] & (~hit)) | (cache_line[k][1934] & (hit));
				cache_line[k][1935] = (mem_line[line_addr][1935] & (~hit)) | (cache_line[k][1935] & (hit));
				cache_line[k][1936] = (mem_line[line_addr][1936] & (~hit)) | (cache_line[k][1936] & (hit));
				cache_line[k][1937] = (mem_line[line_addr][1937] & (~hit)) | (cache_line[k][1937] & (hit));
				cache_line[k][1938] = (mem_line[line_addr][1938] & (~hit)) | (cache_line[k][1938] & (hit));
				cache_line[k][1939] = (mem_line[line_addr][1939] & (~hit)) | (cache_line[k][1939] & (hit));
				cache_line[k][1940] = (mem_line[line_addr][1940] & (~hit)) | (cache_line[k][1940] & (hit));
				cache_line[k][1941] = (mem_line[line_addr][1941] & (~hit)) | (cache_line[k][1941] & (hit));
				cache_line[k][1942] = (mem_line[line_addr][1942] & (~hit)) | (cache_line[k][1942] & (hit));
				cache_line[k][1943] = (mem_line[line_addr][1943] & (~hit)) | (cache_line[k][1943] & (hit));
				cache_line[k][1944] = (mem_line[line_addr][1944] & (~hit)) | (cache_line[k][1944] & (hit));
				cache_line[k][1945] = (mem_line[line_addr][1945] & (~hit)) | (cache_line[k][1945] & (hit));
				cache_line[k][1946] = (mem_line[line_addr][1946] & (~hit)) | (cache_line[k][1946] & (hit));
				cache_line[k][1947] = (mem_line[line_addr][1947] & (~hit)) | (cache_line[k][1947] & (hit));
				cache_line[k][1948] = (mem_line[line_addr][1948] & (~hit)) | (cache_line[k][1948] & (hit));
				cache_line[k][1949] = (mem_line[line_addr][1949] & (~hit)) | (cache_line[k][1949] & (hit));
				cache_line[k][1950] = (mem_line[line_addr][1950] & (~hit)) | (cache_line[k][1950] & (hit));
				cache_line[k][1951] = (mem_line[line_addr][1951] & (~hit)) | (cache_line[k][1951] & (hit));
				cache_line[k][1952] = (mem_line[line_addr][1952] & (~hit)) | (cache_line[k][1952] & (hit));
				cache_line[k][1953] = (mem_line[line_addr][1953] & (~hit)) | (cache_line[k][1953] & (hit));
				cache_line[k][1954] = (mem_line[line_addr][1954] & (~hit)) | (cache_line[k][1954] & (hit));
				cache_line[k][1955] = (mem_line[line_addr][1955] & (~hit)) | (cache_line[k][1955] & (hit));
				cache_line[k][1956] = (mem_line[line_addr][1956] & (~hit)) | (cache_line[k][1956] & (hit));
				cache_line[k][1957] = (mem_line[line_addr][1957] & (~hit)) | (cache_line[k][1957] & (hit));
				cache_line[k][1958] = (mem_line[line_addr][1958] & (~hit)) | (cache_line[k][1958] & (hit));
				cache_line[k][1959] = (mem_line[line_addr][1959] & (~hit)) | (cache_line[k][1959] & (hit));
				cache_line[k][1960] = (mem_line[line_addr][1960] & (~hit)) | (cache_line[k][1960] & (hit));
				cache_line[k][1961] = (mem_line[line_addr][1961] & (~hit)) | (cache_line[k][1961] & (hit));
				cache_line[k][1962] = (mem_line[line_addr][1962] & (~hit)) | (cache_line[k][1962] & (hit));
				cache_line[k][1963] = (mem_line[line_addr][1963] & (~hit)) | (cache_line[k][1963] & (hit));
				cache_line[k][1964] = (mem_line[line_addr][1964] & (~hit)) | (cache_line[k][1964] & (hit));
				cache_line[k][1965] = (mem_line[line_addr][1965] & (~hit)) | (cache_line[k][1965] & (hit));
				cache_line[k][1966] = (mem_line[line_addr][1966] & (~hit)) | (cache_line[k][1966] & (hit));
				cache_line[k][1967] = (mem_line[line_addr][1967] & (~hit)) | (cache_line[k][1967] & (hit));
				cache_line[k][1968] = (mem_line[line_addr][1968] & (~hit)) | (cache_line[k][1968] & (hit));
				cache_line[k][1969] = (mem_line[line_addr][1969] & (~hit)) | (cache_line[k][1969] & (hit));
				cache_line[k][1970] = (mem_line[line_addr][1970] & (~hit)) | (cache_line[k][1970] & (hit));
				cache_line[k][1971] = (mem_line[line_addr][1971] & (~hit)) | (cache_line[k][1971] & (hit));
				cache_line[k][1972] = (mem_line[line_addr][1972] & (~hit)) | (cache_line[k][1972] & (hit));
				cache_line[k][1973] = (mem_line[line_addr][1973] & (~hit)) | (cache_line[k][1973] & (hit));
				cache_line[k][1974] = (mem_line[line_addr][1974] & (~hit)) | (cache_line[k][1974] & (hit));
				cache_line[k][1975] = (mem_line[line_addr][1975] & (~hit)) | (cache_line[k][1975] & (hit));
				cache_line[k][1976] = (mem_line[line_addr][1976] & (~hit)) | (cache_line[k][1976] & (hit));
				cache_line[k][1977] = (mem_line[line_addr][1977] & (~hit)) | (cache_line[k][1977] & (hit));
				cache_line[k][1978] = (mem_line[line_addr][1978] & (~hit)) | (cache_line[k][1978] & (hit));
				cache_line[k][1979] = (mem_line[line_addr][1979] & (~hit)) | (cache_line[k][1979] & (hit));
				cache_line[k][1980] = (mem_line[line_addr][1980] & (~hit)) | (cache_line[k][1980] & (hit));
				cache_line[k][1981] = (mem_line[line_addr][1981] & (~hit)) | (cache_line[k][1981] & (hit));
				cache_line[k][1982] = (mem_line[line_addr][1982] & (~hit)) | (cache_line[k][1982] & (hit));
				cache_line[k][1983] = (mem_line[line_addr][1983] & (~hit)) | (cache_line[k][1983] & (hit));
				cache_line[k][1984] = (mem_line[line_addr][1984] & (~hit)) | (cache_line[k][1984] & (hit));
				cache_line[k][1985] = (mem_line[line_addr][1985] & (~hit)) | (cache_line[k][1985] & (hit));
				cache_line[k][1986] = (mem_line[line_addr][1986] & (~hit)) | (cache_line[k][1986] & (hit));
				cache_line[k][1987] = (mem_line[line_addr][1987] & (~hit)) | (cache_line[k][1987] & (hit));
				cache_line[k][1988] = (mem_line[line_addr][1988] & (~hit)) | (cache_line[k][1988] & (hit));
				cache_line[k][1989] = (mem_line[line_addr][1989] & (~hit)) | (cache_line[k][1989] & (hit));
				cache_line[k][1990] = (mem_line[line_addr][1990] & (~hit)) | (cache_line[k][1990] & (hit));
				cache_line[k][1991] = (mem_line[line_addr][1991] & (~hit)) | (cache_line[k][1991] & (hit));
				cache_line[k][1992] = (mem_line[line_addr][1992] & (~hit)) | (cache_line[k][1992] & (hit));
				cache_line[k][1993] = (mem_line[line_addr][1993] & (~hit)) | (cache_line[k][1993] & (hit));
				cache_line[k][1994] = (mem_line[line_addr][1994] & (~hit)) | (cache_line[k][1994] & (hit));
				cache_line[k][1995] = (mem_line[line_addr][1995] & (~hit)) | (cache_line[k][1995] & (hit));
				cache_line[k][1996] = (mem_line[line_addr][1996] & (~hit)) | (cache_line[k][1996] & (hit));
				cache_line[k][1997] = (mem_line[line_addr][1997] & (~hit)) | (cache_line[k][1997] & (hit));
				cache_line[k][1998] = (mem_line[line_addr][1998] & (~hit)) | (cache_line[k][1998] & (hit));
				cache_line[k][1999] = (mem_line[line_addr][1999] & (~hit)) | (cache_line[k][1999] & (hit));
				cache_line[k][2000] = (mem_line[line_addr][2000] & (~hit)) | (cache_line[k][2000] & (hit));
				cache_line[k][2001] = (mem_line[line_addr][2001] & (~hit)) | (cache_line[k][2001] & (hit));
				cache_line[k][2002] = (mem_line[line_addr][2002] & (~hit)) | (cache_line[k][2002] & (hit));
				cache_line[k][2003] = (mem_line[line_addr][2003] & (~hit)) | (cache_line[k][2003] & (hit));
				cache_line[k][2004] = (mem_line[line_addr][2004] & (~hit)) | (cache_line[k][2004] & (hit));
				cache_line[k][2005] = (mem_line[line_addr][2005] & (~hit)) | (cache_line[k][2005] & (hit));
				cache_line[k][2006] = (mem_line[line_addr][2006] & (~hit)) | (cache_line[k][2006] & (hit));
				cache_line[k][2007] = (mem_line[line_addr][2007] & (~hit)) | (cache_line[k][2007] & (hit));
				cache_line[k][2008] = (mem_line[line_addr][2008] & (~hit)) | (cache_line[k][2008] & (hit));
				cache_line[k][2009] = (mem_line[line_addr][2009] & (~hit)) | (cache_line[k][2009] & (hit));
				cache_line[k][2010] = (mem_line[line_addr][2010] & (~hit)) | (cache_line[k][2010] & (hit));
				cache_line[k][2011] = (mem_line[line_addr][2011] & (~hit)) | (cache_line[k][2011] & (hit));
				cache_line[k][2012] = (mem_line[line_addr][2012] & (~hit)) | (cache_line[k][2012] & (hit));
				cache_line[k][2013] = (mem_line[line_addr][2013] & (~hit)) | (cache_line[k][2013] & (hit));
				cache_line[k][2014] = (mem_line[line_addr][2014] & (~hit)) | (cache_line[k][2014] & (hit));
				cache_line[k][2015] = (mem_line[line_addr][2015] & (~hit)) | (cache_line[k][2015] & (hit));
				cache_line[k][2016] = (mem_line[line_addr][2016] & (~hit)) | (cache_line[k][2016] & (hit));
				cache_line[k][2017] = (mem_line[line_addr][2017] & (~hit)) | (cache_line[k][2017] & (hit));
				cache_line[k][2018] = (mem_line[line_addr][2018] & (~hit)) | (cache_line[k][2018] & (hit));
				cache_line[k][2019] = (mem_line[line_addr][2019] & (~hit)) | (cache_line[k][2019] & (hit));
				cache_line[k][2020] = (mem_line[line_addr][2020] & (~hit)) | (cache_line[k][2020] & (hit));
				cache_line[k][2021] = (mem_line[line_addr][2021] & (~hit)) | (cache_line[k][2021] & (hit));
				cache_line[k][2022] = (mem_line[line_addr][2022] & (~hit)) | (cache_line[k][2022] & (hit));
				cache_line[k][2023] = (mem_line[line_addr][2023] & (~hit)) | (cache_line[k][2023] & (hit));
				cache_line[k][2024] = (mem_line[line_addr][2024] & (~hit)) | (cache_line[k][2024] & (hit));
				cache_line[k][2025] = (mem_line[line_addr][2025] & (~hit)) | (cache_line[k][2025] & (hit));
				cache_line[k][2026] = (mem_line[line_addr][2026] & (~hit)) | (cache_line[k][2026] & (hit));
				cache_line[k][2027] = (mem_line[line_addr][2027] & (~hit)) | (cache_line[k][2027] & (hit));
				cache_line[k][2028] = (mem_line[line_addr][2028] & (~hit)) | (cache_line[k][2028] & (hit));
				cache_line[k][2029] = (mem_line[line_addr][2029] & (~hit)) | (cache_line[k][2029] & (hit));
				cache_line[k][2030] = (mem_line[line_addr][2030] & (~hit)) | (cache_line[k][2030] & (hit));
				cache_line[k][2031] = (mem_line[line_addr][2031] & (~hit)) | (cache_line[k][2031] & (hit));
				cache_line[k][2032] = (mem_line[line_addr][2032] & (~hit)) | (cache_line[k][2032] & (hit));
				cache_line[k][2033] = (mem_line[line_addr][2033] & (~hit)) | (cache_line[k][2033] & (hit));
				cache_line[k][2034] = (mem_line[line_addr][2034] & (~hit)) | (cache_line[k][2034] & (hit));
				cache_line[k][2035] = (mem_line[line_addr][2035] & (~hit)) | (cache_line[k][2035] & (hit));
				cache_line[k][2036] = (mem_line[line_addr][2036] & (~hit)) | (cache_line[k][2036] & (hit));
				cache_line[k][2037] = (mem_line[line_addr][2037] & (~hit)) | (cache_line[k][2037] & (hit));
				cache_line[k][2038] = (mem_line[line_addr][2038] & (~hit)) | (cache_line[k][2038] & (hit));
				cache_line[k][2039] = (mem_line[line_addr][2039] & (~hit)) | (cache_line[k][2039] & (hit));
				cache_line[k][2040] = (mem_line[line_addr][2040] & (~hit)) | (cache_line[k][2040] & (hit));
				cache_line[k][2041] = (mem_line[line_addr][2041] & (~hit)) | (cache_line[k][2041] & (hit));
				cache_line[k][2042] = (mem_line[line_addr][2042] & (~hit)) | (cache_line[k][2042] & (hit));
				cache_line[k][2043] = (mem_line[line_addr][2043] & (~hit)) | (cache_line[k][2043] & (hit));
				cache_line[k][2044] = (mem_line[line_addr][2044] & (~hit)) | (cache_line[k][2044] & (hit));
				cache_line[k][2045] = (mem_line[line_addr][2045] & (~hit)) | (cache_line[k][2045] & (hit));
				cache_line[k][2046] = (mem_line[line_addr][2046] & (~hit)) | (cache_line[k][2046] & (hit));
				cache_line[k][2047] = (mem_line[line_addr][2047] & (~hit)) | (cache_line[k][2047] & (hit));

				tag_array[k] = tag_inp;
				line = cache_line[k];
				//linterest = k;
				//line = mem_line[255];
				//line = cache_line[1];

			//end
	end

	Offset_2_Byte b(line, Block_Offset, ByTe);
	//assign loi = k;

endmodule // direct_cache