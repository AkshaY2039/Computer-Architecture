/*
Computer Architecture Lab 2 - 08-01-2018
	Assignment : Floating Point Adder
	Module : 32b Right Shifter
		-- Eshita Arza	(COE15B013)
		-- Akshay Kumar	(CED15I031)
*/

module right_shifter(x, s, cout, clk);

	input [31:0]x;
	input clk;
	input [4:0]s;
	output [31:0]cout;
	//input enable_right_shift;

	wire [31:0]w1, w2, w3, w4, w5;
	wire [31:0]l1, l2, l3, l4;
	wire [4:0]s1, s2, s3, s4;

	//level 1
	mux m1(x[1], x[0], s[0], w1[0]);
	mux m2(x[2], x[1], s[0], w1[1]);
	mux m3(x[3], x[2], s[0], w1[2]);
	mux m4(x[4], x[3], s[0], w1[3]);
	mux m5(x[5], x[4], s[0], w1[4]);
	mux m6(x[6], x[5], s[0], w1[5]);
	mux m7(x[7], x[6], s[0], w1[6]);
	mux m8(x[8], x[7], s[0], w1[7]);
	mux m9(x[9], x[8], s[0], w1[8]);
	mux m10(x[10], x[9], s[0], w1[9]);
	mux m11(x[11], x[10], s[0], w1[10]);
	mux m12(x[12], x[11], s[0], w1[11]);
	mux m13(x[13], x[12], s[0], w1[12]);
	mux m14(x[14], x[13], s[0], w1[13]);
	mux m15(x[15], x[14], s[0], w1[14]);
	mux m16(x[16], x[15], s[0], w1[15]);
	mux m17(x[17], x[16], s[0], w1[16]);
	mux m18(x[18], x[17], s[0], w1[17]);
	mux m19(x[19], x[18], s[0], w1[18]);
	mux m20(x[20], x[19], s[0], w1[19]);
	mux m21(x[21], x[20], s[0], w1[20]);
	mux m22(x[22], x[21], s[0], w1[21]);
	mux m23(x[23], x[22], s[0], w1[22]);
	mux m24(x[24], x[23], s[0], w1[23]);
	mux m25(x[25], x[24], s[0], w1[24]);
	mux m26(x[26], x[25], s[0], w1[25]);
	mux m27(x[27], x[26], s[0], w1[26]);
	mux m28(x[28], x[27], s[0], w1[27]);
	mux m29(x[29], x[28], s[0], w1[28]);
	mux m30(x[30], x[29], s[0], w1[29]);
	mux m31(x[31], x[30], s[0], w1[30]);
	mux m32(1'b0 , x[31], s[0], w1[31]);

	diff p0(w1[0], l1[0], clk);
	diff p1(w1[1], l1[1], clk);
	diff p2(w1[2], l1[2], clk);
	diff p3(w1[3], l1[3], clk);
	diff p4(w1[4], l1[4], clk);
	diff p5(w1[5], l1[5], clk);
	diff p6(w1[6], l1[6], clk);
	diff p7(w1[7], l1[7], clk);
	diff p8(w1[8], l1[8], clk);
	diff p9(w1[9], l1[9], clk);
	diff p10(w1[10], l1[10], clk);
	diff p11(w1[11], l1[11], clk);
	diff p12(w1[12], l1[12], clk);
	diff p13(w1[13], l1[13], clk);
	diff p14(w1[14], l1[14], clk);
	diff p15(w1[15], l1[15], clk);
	diff p16(w1[16], l1[16], clk);
	diff p17(w1[17], l1[17], clk);
	diff p18(w1[18], l1[18], clk);
	diff p19(w1[19], l1[19], clk);
	diff p20(w1[20], l1[20], clk);
	diff p21(w1[21], l1[21], clk);
	diff p22(w1[22], l1[22], clk);
	diff p23(w1[23], l1[23], clk);
	diff p24(w1[24], l1[24], clk);
	diff p25(w1[25], l1[25], clk);
	diff p26(w1[26], l1[26], clk);
	diff p27(w1[27], l1[27], clk);
	diff p28(w1[28], l1[28], clk);
	diff p29(w1[29], l1[29], clk);
	diff p30(w1[30], l1[30], clk);
	diff p31(w1[31], l1[31], clk);

	diff k1(s[0], s1[0], clk);
	diff k2(s[1], s1[1], clk);
	diff k3(s[2], s1[2], clk);
	diff k4(s[3], s1[3], clk);
	diff k5(s[4], s1[4], clk);

	//level2
	mux mq1(l1[2], l1[0], s1[1], w2[0]);
	mux mq2(l1[3], l1[1], s1[1], w2[1]);
	mux mq3(l1[4], l1[2], s1[1], w2[2]);
	mux mq4(l1[5], l1[3], s1[1], w2[3]);
	mux mq5(l1[6], l1[4], s1[1], w2[4]);
	mux mq6(l1[7], l1[5], s1[1], w2[5]);
	mux mq7(l1[8], l1[6], s1[1], w2[6]);
	mux mq8(l1[9], l1[7], s1[1], w2[7]);
	mux mq9(l1[10], l1[8], s1[1], w2[8]);
	mux mq10(l1[11], l1[9], s1[1], w2[9]);
	mux mq11(l1[12], l1[10], s1[1], w2[10]);
	mux mq12(l1[13], l1[11], s1[1], w2[11]);
	mux mq13(l1[14], l1[12], s1[1], w2[12]);
	mux mq14(l1[15], l1[13], s1[1], w2[13]);
	mux mq15(l1[16], l1[14], s1[1], w2[14]);
	mux mq16(l1[17], l1[15], s1[1], w2[15]);
	mux mq17(l1[18], l1[16], s1[1], w2[16]);
	mux mq18(l1[19], l1[17], s1[1], w2[17]);
	mux mq19(l1[20], l1[18], s1[1], w2[18]);
	mux mq20(l1[21], l1[19], s1[1], w2[19]);
	mux mq21(l1[22], l1[20], s1[1], w2[20]);
	mux mq22(l1[23], l1[21], s1[1], w2[21]);
	mux mq23(l1[24], l1[22], s1[1], w2[22]);
	mux mq24(l1[25], l1[23], s1[1], w2[23]);
	mux mq25(l1[26], l1[24], s1[1], w2[24]);
	mux mq26(l1[27], l1[25], s1[1], w2[25]);
	mux mq27(l1[28], l1[26], s1[1], w2[26]);
	mux mq28(l1[29], l1[27], s1[1], w2[27]);
	mux mq29(l1[30], l1[28], s1[1], w2[28]);
	mux mq30(l1[31], l1[29], s1[1], w2[29]);
	mux mq31(1'b0, l1[30], s1[1], w2[30]);
	mux mq32(1'b0, l1[31], s1[1], w2[31]);

	diff qp0(w2[0], l2[0], clk);
	diff qp1(w2[1], l2[1], clk);
	diff qp2(w2[2], l2[2], clk);
	diff qp3(w2[3], l2[3], clk);
	diff qp4(w2[4], l2[4], clk);
	diff qp5(w2[5], l2[5], clk);
	diff qp6(w2[6], l2[6], clk);
	diff qp7(w2[7], l2[7], clk);
	diff qp8(w2[8], l2[8], clk);
	diff qp9(w2[9], l2[9], clk);
	diff qp10(w2[10], l2[10], clk);
	diff qp11(w2[11], l2[11], clk);
	diff qp12(w2[12], l2[12], clk);
	diff qp13(w2[13], l2[13], clk);
	diff qp14(w2[14], l2[14], clk);
	diff qp15(w2[15], l2[15], clk);
	diff qp16(w2[16], l2[16], clk);
	diff qp17(w2[17], l2[17], clk);
	diff qp18(w2[18], l2[18], clk);
	diff qp19(w2[19], l2[19], clk);
	diff qp20(w2[20], l2[20], clk);
	diff qp21(w2[21], l2[21], clk);
	diff qp22(w2[22], l2[22], clk);
	diff qp23(w2[23], l2[23], clk);
	diff qp24(w2[24], l2[24], clk);
	diff qp25(w2[25], l2[25], clk);
	diff qp26(w2[26], l2[26], clk);
	diff qp27(w2[27], l2[27], clk);
	diff qp28(w2[28], l2[28], clk);
	diff qp29(w2[29], l2[29], clk);
	diff qp30(w2[30], l2[30], clk);
	diff qp31(w2[31], l2[31], clk);

	diff kq1(s1[0], s2[0], clk);
	diff kq2(s1[1], s2[1], clk);
	diff kq3(s1[2], s2[2], clk);
	diff kq4(s1[3], s2[3], clk);
	diff kq5(s1[4], s2[4], clk);

	//level 3
	mux mw1(l2[4], l2[0], s2[2], w3[0]);
	mux mw2(l2[5], l2[1], s2[2], w3[1]);
	mux mw3(l2[6], l2[2], s2[2], w3[2]);
	mux mw4(l2[7], l2[3], s2[2], w3[3]);
	mux mw5(l2[8], l2[4], s2[2], w3[4]);
	mux mw6(l2[9], l2[5], s2[2], w3[5]);
	mux mw7(l2[10], l2[6], s2[2], w3[6]);
	mux mw8(l2[11], l2[7], s2[2], w3[7]);
	mux mw9(l2[12], l2[8], s2[2], w3[8]);
	mux mw10(l2[13], l2[9], s2[2], w3[9]);
	mux mw11(l2[14], l2[10], s2[2], w3[10]);
	mux mw12(l2[15], l2[11], s2[2], w3[11]);
	mux mw13(l2[16], l2[12], s2[2], w3[12]);
	mux mw14(l2[17], l2[13], s2[2], w3[13]);
	mux mw15(l2[18], l2[14], s2[2], w3[14]);
	mux mw16(l2[19], l2[15], s2[2], w3[15]);
	mux mw17(l2[20], l2[16], s2[2], w3[16]);
	mux mw18(l2[21], l2[17], s2[2], w3[17]);
	mux mw19(l2[22], l2[18], s2[2], w3[18]);
	mux mw20(l2[23], l2[19], s2[2], w3[19]);
	mux mw21(l2[24], l2[20], s2[2], w3[20]);
	mux mw22(l2[25], l2[21], s2[2], w3[21]);
	mux mw23(l2[26], l2[22], s2[2], w3[22]);
	mux mw24(l2[27], l2[23], s2[2], w3[23]);
	mux mw25(l2[28], l2[24], s2[2], w3[24]);
	mux mw26(l2[29], l2[25], s2[2], w3[25]);
	mux mw27(l2[30], l2[26], s2[2], w3[26]);
	mux mw28(l2[31], l2[27], s2[2], w3[27]);
	mux mw29(1'b0, l2[28], s2[2], w3[28]);
	mux mw30(1'b0, l2[29], s2[2], w3[29]);
	mux mw31(1'b0, l2[30], s2[2], w3[30]);
	mux mw32(1'b0, l2[31], s2[2], w3[31]);

	diff bp0(w3[0], l3[0], clk);
	diff bp1(w3[1], l3[1], clk);
	diff bp2(w3[2], l3[2], clk);
	diff bp3(w3[3], l3[3], clk);
	diff bp4(w3[4], l3[4], clk);
	diff bp5(w3[5], l3[5], clk);
	diff bp6(w3[6], l3[6], clk);
	diff bp7(w3[7], l3[7], clk);
	diff bp8(w3[8], l3[8], clk);
	diff bp9(w3[9], l3[9], clk);
	diff bp10(w3[10], l3[10], clk);
	diff bp11(w3[11], l3[11], clk);
	diff bp12(w3[12], l3[12], clk);
	diff bp13(w3[13], l3[13], clk);
	diff bp14(w3[14], l3[14], clk);
	diff bp15(w3[15], l3[15], clk);
	diff bp16(w3[16], l3[16], clk);
	diff bp17(w3[17], l3[17], clk);
	diff bp18(w3[18], l3[18], clk);
	diff bp19(w3[19], l3[19], clk);
	diff bp20(w3[20], l3[20], clk);
	diff bp21(w3[21], l3[21], clk);
	diff bp22(w3[22], l3[22], clk);
	diff bp23(w3[23], l3[23], clk);
	diff bp24(w3[24], l3[24], clk);
	diff bp25(w3[25], l3[25], clk);
	diff bp26(w3[26], l3[26], clk);
	diff bp27(w3[27], l3[27], clk);
	diff bp28(w3[28], l3[28], clk);
	diff bp29(w3[29], l3[29], clk);
	diff bp30(w3[30], l3[30], clk);
	diff bp31(w3[31], l3[31], clk);

	diff zq1(s2[0], s3[0], clk);
	diff zq2(s2[1], s3[1], clk);
	diff zq3(s2[2], s3[2], clk);
	diff zq4(s2[3], s3[3], clk);
	diff zq5(s2[4], s3[4], clk);

	//level 4
	mux mr1(l3[8], l3[0], s3[3], w4[0]);
	mux mr2(l3[9], l3[1], s3[3], w4[1]);
	mux mr3(l3[10], l3[2], s3[3], w4[2]);
	mux mr4(l3[11], l3[3], s3[3], w4[3]);
	mux mr5(l3[12], l3[4], s3[3], w4[4]);
	mux mr6(l3[13], l3[5], s3[3], w4[5]);
	mux mr7(l3[14], l3[6], s3[3], w4[6]);
	mux mr8(l3[15], l3[7], s3[3], w4[7]);
	mux mr9(l3[16], l3[8], s3[3], w4[8]);
	mux mr10(l3[17], l3[9], s3[3], w4[9]);
	mux mr11(l3[18], l3[10], s3[3], w4[10]);
	mux mr12(l3[19], l3[11], s3[3], w4[11]);
	mux mr13(l3[20], l3[12], s3[3], w4[12]);
	mux mr14(l3[21], l3[13], s3[3], w4[13]);
	mux mr15(l3[22], l3[14], s3[3], w4[14]);
	mux mr16(l3[23], l3[15], s3[3], w4[15]);
	mux mr17(l3[24], l3[16], s3[3], w4[16]);
	mux mr18(l3[25], l3[17], s3[3], w4[17]);
	mux mr19(l3[26], l3[18], s3[3], w4[18]);
	mux mr20(l3[27], l3[19], s3[3], w4[19]);
	mux mr21(l3[28], l3[20], s3[3], w4[20]);
	mux mr22(l3[29], l3[21], s3[3], w4[21]);
	mux mr23(l3[30], l3[22], s3[3], w4[22]);
	mux mr24(l3[31], l3[23], s3[3], w4[23]);
	mux mr25(1'b0, l3[24], s3[3], w4[24]);
	mux mr26(1'b0, l3[25], s3[3], w4[25]);
	mux mr27(1'b0, l3[26], s3[3], w4[26]);
	mux mr28(1'b0, l3[27], s3[3], w4[27]);
	mux mr29(1'b0, l3[28], s3[3], w4[28]);
	mux mr30(1'b0, l3[29], s3[3], w4[29]);
	mux mr31(1'b0, l3[30], s3[3], w4[30]);
	mux mr32(1'b0, l3[31], s3[3], w4[31]);

	diff cp0(w4[0], l4[0], clk);
	diff cp1(w4[1], l4[1], clk);
	diff cp2(w4[2], l4[2], clk);
	diff cp3(w4[3], l4[3], clk);
	diff cp4(w4[4], l4[4], clk);
	diff cp5(w4[5], l4[5], clk);
	diff cp6(w4[6], l4[6], clk);
	diff cp7(w4[7], l4[7], clk);
	diff cp8(w4[8], l4[8], clk);
	diff cp9(w4[9], l4[9], clk);
	diff cp10(w4[10], l4[10], clk);
	diff cp11(w4[11], l4[11], clk);
	diff cp12(w4[12], l4[12], clk);
	diff cp13(w4[13], l4[13], clk);
	diff cp14(w4[14], l4[14], clk);
	diff cp15(w4[15], l4[15], clk);
	diff cp16(w4[16], l4[16], clk);
	diff cp17(w4[17], l4[17], clk);
	diff cp18(w4[18], l4[18], clk);
	diff cp19(w4[19], l4[19], clk);
	diff cp20(w4[20], l4[20], clk);
	diff cp21(w4[21], l4[21], clk);
	diff cp22(w4[22], l4[22], clk);
	diff cp23(w4[23], l4[23], clk);
	diff cp24(w4[24], l4[24], clk);
	diff cp25(w4[25], l4[25], clk);
	diff cp26(w4[26], l4[26], clk);
	diff cp27(w4[27], l4[27], clk);
	diff cp28(w4[28], l4[28], clk);
	diff cp29(w4[29], l4[29], clk);
	diff cp30(w4[30], l4[30], clk);
	diff cp31(w4[31], l4[31], clk);

	diff xq1(s3[0], s4[0], clk);
	diff xq2(s3[1], s4[1], clk);
	diff xq3(s3[2], s4[2], clk);
	diff xq4(s3[3], s4[3], clk);
	diff xq5(s3[4], s4[4], clk);

	//level 5
	mux mp1(l4[16], l4[0], s4[4], w5[0]);
	mux mp2(l4[17], l4[1], s4[4], w5[1]);
	mux mp3(l4[18], l4[2], s4[4], w5[2]);
	mux mp4(l4[19], l4[3], s4[4], w5[3]);
	mux mp5(l4[20], l4[4], s4[4], w5[4]);
	mux mp6(l4[21], l4[5], s4[4], w5[5]);
	mux mp7(l4[22], l4[6], s4[4], w5[6]);
	mux mp8(l4[23], l4[7], s4[4], w5[7]);
	mux mp9(l4[24], l4[8], s4[4], w5[8]);
	mux mp10(l4[25], l4[9], s4[4], w5[9]);
	mux mp11(l4[26], l4[10], s4[4], w5[10]);
	mux mp12(l4[27], l4[11], s4[4], w5[11]);
	mux mp13(l4[28], l4[12], s4[4], w5[12]);
	mux mp14(l4[28], l4[13], s4[4], w5[13]);
	mux mp15(l4[29], l4[14], s4[4], w5[14]);
	mux mp16(l4[30], l4[15], s4[4], w5[15]);
	mux mp17(l4[31], l4[16], s4[4], w5[16]);
	mux mp18(1'b0, l4[17], s4[4], w5[17]);
	mux mp19(1'b0, l4[18], s4[4], w5[18]);
	mux mp20(1'b0, l4[19], s4[4], w5[19]);
	mux mp21(1'b0, l4[20], s4[4], w5[20]);
	mux mp22(1'b0, l4[21], s4[4], w5[21]);
	mux mp23(1'b0, l4[22], s4[4], w5[22]);
	mux mp24(1'b0, l4[23], s4[4], w5[23]);
	mux mp25(1'b0, l4[24], s4[4], w5[24]);
	mux mp26(1'b0, l4[25], s4[4], w5[25]);
	mux mp27(1'b0, l4[26], s4[4], w5[26]);
	mux mp28(1'b0, l4[27], s4[4], w5[27]);
	mux mp29(1'b0, l4[28], s4[4], w5[28]);
	mux mp30(1'b0, l4[29], s4[4], w5[29]);
	mux mp31(1'b0, l4[30], s4[4], w5[30]);
	mux mp32(1'b0, l4[31], s4[4], w5[31]);

	assign cout = w5;

endmodule // right_shifter