/*
Computer Architecture Lab 2 - 08-01-2018
	Assignment : Floating Point Multiplier
	Module : 64b Carry Save Adder
		-- Eshita Arza	(COE15B013)
		-- Akshay Kumar	(CED15I031)
*/

module csa(x, y, z, s, c);

	input [63:0]x, y, z;
	input cin;
	output [63:0]s;
	output [64:0]c;

	assign s = x ^ y ^ z;
	assign c[0] = 1'b0;
	assign c[1] = (x[0] & y[0]) | (y[0] & z[0]) | (z[0] & x[0]);
	assign c[2] = (x[1] & y[1]) | (y[1] & z[1]) | (z[1] & x[1]);
	assign c[3] = (x[2] & y[2]) | (y[2] & z[2]) | (z[2] & x[2]);
	assign c[4] = (x[3] & y[3]) | (y[3] & z[3]) | (z[3] & x[3]);
	assign c[5] = (x[4] & y[4]) | (y[4] & z[4]) | (z[4] & x[4]);
	assign c[6] = (x[5] & y[5]) | (y[5] & z[5]) | (z[5] & x[5]);
	assign c[7] = (x[6] & y[6]) | (y[6] & z[6]) | (z[6] & x[6]);
	assign c[8] = (x[7] & y[7]) | (y[7] & z[7]) | (z[7] & x[7]);
	assign c[9] = (x[8] & y[8]) | (y[8] & z[8]) | (z[8] & x[8]);
	assign c[10] = (x[9] & y[9]) | (y[9] & z[9]) | (z[9] & x[9]);
	assign c[11] = (x[10] & y[10]) | (y[10] & z[10]) | (z[10] & x[10]);
	assign c[12] = (x[11] & y[11]) | (y[11] & z[11]) | (z[11] & x[11]);
	assign c[13] = (x[12] & y[12]) | (y[12] & z[12]) | (z[12] & x[12]);
	assign c[14] = (x[13] & y[13]) | (y[13] & z[13]) | (z[13] & x[13]);
	assign c[15] = (x[14] & y[14]) | (y[14] & z[14]) | (z[14] & x[14]);
	assign c[16] = (x[15] & y[15]) | (y[15] & z[15]) | (z[15] & x[15]);
	assign c[17] = (x[16] & y[16]) | (y[16] & z[16]) | (z[16] & x[16]);
	assign c[18] = (x[17] & y[17]) | (y[17] & z[17]) | (z[17] & x[17]);
	assign c[19] = (x[18] & y[18]) | (y[18] & z[18]) | (z[18] & x[18]);
	assign c[20] = (x[19] & y[19]) | (y[19] & z[19]) | (z[19] & x[19]);
	assign c[21] = (x[20] & y[20]) | (y[20] & z[20]) | (z[20] & x[20]);
	assign c[22] = (x[21] & y[21]) | (y[21] & z[21]) | (z[21] & x[21]);
	assign c[23] = (x[22] & y[22]) | (y[22] & z[22]) | (z[22] & x[22]);
	assign c[24] = (x[23] & y[23]) | (y[23] & z[23]) | (z[23] & x[23]);
	assign c[25] = (x[24] & y[24]) | (y[24] & z[24]) | (z[24] & x[24]);
	assign c[26] = (x[25] & y[25]) | (y[25] & z[25]) | (z[25] & x[25]);
	assign c[27] = (x[26] & y[26]) | (y[26] & z[26]) | (z[26] & x[26]);
	assign c[28] = (x[27] & y[27]) | (y[27] & z[27]) | (z[27] & x[27]);
	assign c[29] = (x[28] & y[28]) | (y[28] & z[28]) | (z[28] & x[28]);
	assign c[30] = (x[29] & y[29]) | (y[29] & z[29]) | (z[29] & x[29]);
	assign c[31] = (x[30] & y[30]) | (y[30] & z[30]) | (z[30] & x[30]);
	assign c[32] = (x[31] & y[31]) | (y[31] & z[31]) | (z[31] & x[31]);
	assign c[33] = (x[32] & y[32]) | (y[32] & z[32]) | (z[32] & x[32]);
	assign c[34] = (x[33] & y[33]) | (y[33] & z[33]) | (z[33] & x[33]);
	assign c[35] = (x[34] & y[34]) | (y[34] & z[34]) | (z[34] & x[34]);
	assign c[36] = (x[35] & y[35]) | (y[35] & z[35]) | (z[35] & x[35]);
	assign c[37] = (x[36] & y[36]) | (y[36] & z[36]) | (z[36] & x[36]);
	assign c[38] = (x[37] & y[37]) | (y[37] & z[37]) | (z[37] & x[37]);
	assign c[39] = (x[38] & y[38]) | (y[38] & z[38]) | (z[38] & x[38]);
	assign c[40] = (x[39] & y[39]) | (y[39] & z[39]) | (z[39] & x[39]);
	assign c[41] = (x[40] & y[40]) | (y[40] & z[40]) | (z[40] & x[40]);
	assign c[42] = (x[41] & y[41]) | (y[41] & z[41]) | (z[41] & x[41]);
	assign c[43] = (x[42] & y[42]) | (y[42] & z[42]) | (z[42] & x[42]);
	assign c[44] = (x[43] & y[43]) | (y[43] & z[43]) | (z[43] & x[43]);
	assign c[45] = (x[44] & y[44]) | (y[44] & z[44]) | (z[44] & x[44]);
	assign c[46] = (x[45] & y[45]) | (y[45] & z[45]) | (z[45] & x[45]);
	assign c[47] = (x[46] & y[46]) | (y[46] & z[46]) | (z[46] & x[46]);
	assign c[48] = (x[47] & y[47]) | (y[47] & z[47]) | (z[47] & x[47]);
	assign c[49] = (x[48] & y[48]) | (y[48] & z[48]) | (z[48] & x[48]);
	assign c[50] = (x[49] & y[49]) | (y[49] & z[49]) | (z[49] & x[49]);
	assign c[51] = (x[50] & y[50]) | (y[50] & z[50]) | (z[50] & x[50]);
	assign c[52] = (x[51] & y[51]) | (y[51] & z[51]) | (z[51] & x[51]);
	assign c[53] = (x[52] & y[52]) | (y[52] & z[52]) | (z[52] & x[52]);
	assign c[54] = (x[53] & y[53]) | (y[53] & z[53]) | (z[53] & x[53]);
	assign c[55] = (x[54] & y[54]) | (y[54] & z[54]) | (z[54] & x[54]);
	assign c[56] = (x[55] & y[55]) | (y[55] & z[55]) | (z[55] & x[55]);
	assign c[57] = (x[56] & y[56]) | (y[56] & z[56]) | (z[56] & x[56]);
	assign c[58] = (x[57] & y[57]) | (y[57] & z[57]) | (z[57] & x[57]);
	assign c[59] = (x[58] & y[58]) | (y[58] & z[58]) | (z[58] & x[58]);
	assign c[60] = (x[59] & y[59]) | (y[59] & z[59]) | (z[59] & x[59]);
	assign c[61] = (x[60] & y[60]) | (y[60] & z[60]) | (z[60] & x[60]);
	assign c[62] = (x[61] & y[61]) | (y[61] & z[61]) | (z[61] & x[61]);
	assign c[63] = (x[62] & y[62]) | (y[62] & z[62]) | (z[62] & x[62]);
	assign c[64] = (x[63] & y[63]) | (y[63] & z[63]) | (z[63] & x[63]);

endmodule // csa